PK   }Q�TP�d�'  �    cirkitFile.json�]]s�Fr�+)�UPa�0�}���U~HֵNm���fE�n(j���{ )�A6���[�===�����j_��{\7O�n��n��{z\}�n�s�o�/��߭��ׇ��O���ϫO���g�|�;��͓��ZumQ+!���晶Fg�f�gj�V7֪�^��|���׻������!_K6.B�Vl\�|����ڰ9p�u���E�ז́���K6.B�����G�%± �J��|gɆp,���X�&±�L6�c�w�lǂ�6���q�!��dC���w�!��dC8��&�wJ��dC8|�Ɇp,����X�}'±��N6�c���lǂ�;�oO�v�l_�������C�������{�~b�	,;�{k�~����=�m�7u�mV�U�i��Y�k�5ۍ6Ji�H�@��V����]LO��Vm�Q٦������:ϳjc뮭��-���t�����������Xv�Zau�����lL�*���6�R+WY�6�5�����R���I��IL��Ic[Lc[,`7ۏs[�b�ٰj7X�C�	,�|]`uW`ue'������bue'���u��]��������VwVwPvˮ�1 ����O���{`���0R&[7���͔�J7�1e�"�&�,e�i��+f�#���o��U����D���T܅p,&���� �������FX~̯�I��`�	0�~�?p���'"�b���:7�-2�X�i]6Yi�*3f�1�V���u��$����_�e�8T��~1���4���f��L���F�&�J����6ʲ�8��H�OD�E��V���Yc��p��&�ۍ�r][�IY�v���}p�&�a�� ��U���B~�M��Y�}��,	X��M��_tw��]�T6�D�f��*+kYd]k[Y��,�@�V=x�L��4	Ӱ��_��?p���'"�fw����$8���Teڮ�l'2!��L��f[dM���z+�2�W�y�UC~э[kM^�u��*Ӆl�M۔Y��
7W�؆��;hJpp��'���3y`���C,?�7�+�688����OD�� �q�ĳ'���_�ϊO���{����ٓ��\j�}���0�x�.���z���s��^r�VY���<Yp�<ܘ��h�z����[3�~p�m���;S��߆��}fGnoM�~���Nv�.��H�V�G�T_#=�e�2��H�f���.U4��Yg��p�j��O�:�֔��M�Ѫ���dEџ��u��BWY�X����6Uۻ&γֳ�ٖB�T��:P�y��/@M��2��*=	'�y��4��}== }=�_��(�{�2at�[�&+����m%�+�o�3ғS��������.zӔn�f��0�"w>�u:7�4������)�Bz2K������Mɉ_O�pZ�v1f�2٦}?=٦�h��125&QG4γֳӓ|b_e�)��*��)��H�Be)�xm�$�<D��sL85�'TCHMd��3�ɩ(����Pw�yrꝉKX�'�LL�&�#��~VP�<1��t������yt���9��O<q5�����I��NQ�;�4�I���G<�]��Q�������p� h��x�dP�\[�H31�b�AR��<f�H�,�v&�IE�v	iKu���G�� ����<0���%� �
���9CzjE<
�Ԃ!��ۮL�Ir�$*��#���kGĻ�LEx����>p�S�7OO{~j�տ�ÿ��| �#�`�����4DF �!��0��1�@@C�q#А��4$&�0Ӕ�\$�k��6�o��F!��8�|��9o�1�9���G!��8�|��9q�1I:�̏K�G!��8��߸	8̏K�G!S��8�����q�1;�̏K�G!S��8���������V~�8�pA
�&s���r���?�F�~~�B��}E���؀ѫ�|��%����1��1�Q�z�"�5ƕo�~��^�d��\z]�k���
��\����	�@�.�5̌�р�=�
��\ì��Y�@�.�5̨�р�2�
��\�l��2W��,r-�6�����Ba�l#��H�.zE��
�	���� %,�6�g��e� �9H	K���`)a� ,�xR�2a�"l#i��H�.�E���2�X����e±E�Fr��a��]&$����2AY����e²([���2qY����L\��Hv<,R���e����X��"u���v�=� G9��e�E�F��a��]&.���e��eA�q�B���L\d ��"u���v�=� �8��e�E�Fң�a��]&.����e� �8H	��eQ��n�'8�������8}==�9 E�����6J�"��{�2��-Jժe8[��Z]+���[eݕ��z��(^��o��֌��ĩ��0>^�D�7#>���\�V5��\�0Zs`N>ضÁ�Ǯ��<W��0��Z�ъ��������Vf�b��[�b3Xqm��,V��ʊ�R�{3�4#`n�$�9�(.7�j"g �>�Jʩ7՝Mtj��K۲�����(7{92c��g5��}ˑ��_w�����_����zw��$�ޝ�酯,���׃'jZ��3j���.��m�zKS3�^��Yp�OԌ��c'jr���B�+{}�JM{}M��z=6�&n�Ps�^�G����ۈ���"n����g��d�׵K�z�cSx^�s��8o�]b"��V��7�b:��p�L��߈�D�rs�����g fa���y(���[&��C}� ���þ~��7/" �8�A���c'��8C���c:��8?�03!B����!�@@�L�F �c&D#�)"�E�6�m����9n�)"��w��F!�2!b8����9p�)"�̇�G!�2!b8�����q�)"�n���������q�)"�̏K�G!�2!b8�����q�)"�̏K�O!2!�Q��"��L�hT�H&D4*P�Kp�dB�h �J�F�u	��L�רШ@�.�5�	���
��%�F2!B4\�B����H&D���ShT�^��Ʉ�@pm
�
��\#�!�L�Q�z]�k$"D�u)4*P�Kp�dB����	��܂�9�2!�"lc��H�.v-w���H�.z-�6�	���2��"lc��H�.�-�6�	���2a�"lc��H�.�-�6�	���2��"lc��H�.�-�6�	���2a�"lc��ȝ�e�E��2!�a��]&.[�m,"�ۅ�Ė���܂pX�n���a˄�E�v��l��L�pX�n���a˄�E�v��l��L�pX�n���a˄�E�v��l��L�pX�n���HlgdB�$�r�Ȅ�GI����	���8�<#"%q�wF&D>J�l�L� ���.��Ʉ��p�vԜL� ����Ʉ�z+Nݧ��	 ����E�9�0+N����	 ��b��buӊə�(.7;9"�fw"gB���L�L�|��]��	`u ��X��Y=" c��g5�L�Waș�(7���	����r��ș�(7߈�	����rS��L�WQș�(7�B΄�G��妷#gB��B΄�G�m��L�|���B΄�G��w����䩙�(��Zj&ī(�L�|��oD΄x�3P3!�Qn�]j&D>ʥ�������úyzxگw��W���[���w��ouӵ����i�v�էϟSND��n��+�L<�8����<����y2�&���`:`g,H0!�c�f����HP!u��[���+RVK�A��q�pH��8�Q���,��Vh�����z1��Q)HT�A$���1a*E�|-mLg1�i��6�a1�$��,ޡu�����]Σ%��2g=�3;f>��֢d=�U
����Z�M�8���q�̉��ԓ�;@�s �g�JL&ߛ�p�:�����
�r��y�'��q�I�K��/#�ٲN�p�"֣��:���!�ԸE[��M�iq�GŻ���y�u������]׏ml���#턇��,� s%�*��X�0�F�i���l�=������&��oP8<Yu� �l���>dٜ��z~�ч,����ү�G,���W֯2��v>#�:�UF��~]G��~��G,��	�����X���ȧ�f�^7�j�S 6�|�}����0��ǶB���g�����-�]���cs�O���q���lu (pw<��C��>����`n��	pwC�k�M~���Ƿ�-~���)�>2~Ć	�|ߤ�9������i�|������O���q����e׮>�����������K����!����,��{_Ll��1&6�����xo�ɂ��ԙ,��p͝ɂ���,��p͞ɂ���s��{"�'�
��c��L\ * N���spy �� 8R>F~�!����L��1����J�?�c�*�sy 棈	)��J�?�c���sy ���S>ƩJ=���J�?�c���sy ����czj۠|�{���4��;��G��ԁ��A�
�:�R����_?����ݜ�
)9��nP���],�H�y��u)px���Ή=����D
�3���`j7�罾��C�5(F�Ã��/RE���A�	DX~�j����J�� ���T�g�oP8���_��;�}��8<����"U޹Sgth�J�N����a��;���b���c�ہ���Ø���Fܠׄй�2��h�2:z	+�s_�0V�����%�h�}et�f����������j�-�ʀ�J�s_̈́�ɹ���gB��Y�֊c5Թ*EG8`����JY7Ac�ӹ���0V(����',7�}�!����G�<a�q  F�Co���cT�y���\��C0�X�s  F��'d��y�� :
k�s50�4�\/��9bT0�T��X�U7bT���cÚ�����g��ḛ8W���0V��S)�nsp�w�P���S������[���ɹS����)����,��+���ȒW�p���p��s�v����.Ks�;�;3 8�= 8]=�k�����iD�cYIhł�)dhł�+dhŒ��A�x��&*��\�p�I?$C.��;<Θ0��ޗ�a�P�l)����C:wN��LJ�%�9��>�ʸA.p>nќ��'�`9/�P���\�܃K�/�:G�����߿�{�%�Y \�6�8g��r���4N/v�xAr�sZ"�;�u!r�s�]$ؑ+�{p��\
�CK��k�Ӝ#�8���p��*���&��r�\b�J����IBw���vG���l�)�%�=v	ݑk�{��#Y��%�\m݃K8`r�u.����=�� b��"А+�{�"�����˦:�F��*XA-��lj��Vm��	3&�o��R�9������ȍZ��c�
����=��$�\�݃K�1�ֻ���ݑ��{�R�Z��cǁ�2'��|?T�׀�ٵ}�<����ͣ��O�W���[�������멷��t���w��C~ep��0>x�a�ԇe�a���a���a67L��I�0�f�S�?äe�j���׊2i��wϤL�ߞ�@�܎I�/Q朣�P&Z�*��p{O��P��1U�p(����/Q�g�%�
�D�����r쑏ݡ�k'��<74��@����2�a� ���r�C\4) ��>��R��pء�)��)���v�"K�2�)>��R���C_�ى�8�!��v���C�2�R#Ňh
إ��)��K�Q�) �t�P3) ���P?) �d?�tQ@.5N�K��Mj\x�r>>�ޥ�O�&��ߥ�O��pK�lR~�=��dRn�=JdR��}�tR����
�ƍw)�I���(�I���(#�Q��{�
ؤ<�
ؤ<�
�$cޣ�P�&�ߥQ�&9��rD��k���Do+�����C��������������/�r�O��#~$O��#u�H���G:�Ȝ>2�G��"�Ȟ>��G��2��:}T��6D��P�*D�"B���FD�q~o��8���\�U)B]��VD�qV��"�z��^�Y/2ԋ|��P/��E��"C��������Yg2ԙ<�L�:�g��P/��E���B���^T�u֋
��^;P�u֋
���zQ�^�Y/�M���a}��|��}Z?����V�m'ݐ+�͑.�j[n3�ɷBئ�u�.�Z��k�ҹ���C�=��DGՇu�o��^W��Z��_��9��%��꿟�Tj��߆?������nؗ���c���i;?��ǟ�.�_���O�V�^����9^w�������ӯ~�7������;��s����y�y�^�����e���է�{�|�ԏ/ۺ9�����_����C[o�/�ÿ|�ؾ��q/�g�h�1qw�=9}|.����1�0��	s�ieg]��i�'��CX���ʷ]�U�γ�uCUvu�4���Q��Q�=>���������ɽ��>[�L��훇�Ԭ�m�C%�w��B���yu���A�v�/�������%��}��,���?fBT��'0��������n� J#�\�<�-�I���,�:{)qi�*d�܏��[���ٓ��f�(r[���o��I�|����`��A����b�]�u���u�<��s���ڽ��_�.u���e�ɚ��L7��6����P�V���.H�%�p_�_Y�o?���ª��S߉��(*UIs��=�BJ��;)�K�"9m΃�1"7�/�e��u߰��GR�%�Ϋ�K7]I���f�>,���	��{�v��!���J�de���؋K�mu+�����8?��ˬQz��^$T�L}���nI�t(}8?vU�{���n�;d�"��,n0荵(�l�X�n'���{k�&���r4�*/�E�vc��S�u�����?��Q�/�X��o-�c�$/��A\N���$E�t�C,U2�b����,Ӑ15SR1eE�,�O�Ӑ1S�-�,I���i�DACE�TDIEDDUUIE,�����߸�;*��`���+�F�<.��`��C����?����x���?}�����>6���<�{�����sS��AѶ]S�f��uV�(Wl�����J�nL�H��	���������o�p���U.�����~*/+yo��l~zm�Amq/�u�yS����	�&�tyo�J�>T�	�������8�����Х<G06!gM�J��/�'�Pr�N�Dg�u/U����U/&��UO.j��){�R�jʝ%]���>��g�.~:��)����׀{'Q8u�=���:���˹�� �����G<��z :��ȫ�r��ZHѯ7�"�*[ݻ��4�0e��j��DSf��n�ۺ�Ô�9b�mL�ltt1�%J�"�!J�ڛH�f��!O~$���)H�Z���p����U�V���|��7��F�6E�t[�<��gV4��L'����ܺ -�	�hwEy\�qz��?������K��8��$��/*��]3��VF�ظ�ʶ����8���6����i�*��t���j	)6�g-w.��__��_��|T�t�/w�!����N/4ъ��l�Y���1��Y�L��Jm�3[� �ܗ�5����sh$U1؈�M�R^�9��_!�>k"���yw|���H�Dڧ_�&$b�L��������~D�r����/"ӕ�S�f�.tv]�)%W��0Ƿ�Lr��J5n�m\���ԙ��L�����
��H7�l��7���W�a�u�c�(zwh��kXq����rXW���{��Ӿ~<5��⫛����:�S�r��dWu�jMf��8��|�׉;7�����<H�I�A?���n���0a�|���$�����ӽ���?��,�d]+8�Q���κqх�uO��VD��ܶ"�*�^Z�X7ֵ:k��݀P���G��F�{���ŝ��8�R곷����M�g��y��tU�~��(���"n[�%����Fvxr�ʌJ7.��bCp+������=�<��}�"�^?wà耝�|������c����v��ܵ|ݗ�a�������]�c�o_\�xx�Y}����������⌰�~�=~�;�9�u��U(���j_��#����w�oO�������/_���c�����б���~����":vz_{r/q���K'�����5$��2��b�r_���_V�;���s��)��	��)���Y�6Z�I�/f�X���a�RD���	�A��}�4���2�j�T l'��P�.�u��b�X��L�b&�LyC*���Q�!�K�c����̖k�*j��s�T��L�bF��&��+-/�\�4t{��h�1�֎���4�/UE��h��(E5�IC.-i�t��1wW��D�N5���k��I�I�4	�7�!IY��z�5iR����(X3,gz�	\�f�;��Q��mn_*n�U.	�Г�2����-MjoHK��5�b�7��i��S�P��P��P��p,eu��Uv��N��I���f(��t�H3�Н�ϡ�����&�r�fH-���Qa�G�^�\���;�xF�&i<r�y�b*���xRG�Zd��%���ܕ�	\�6�X��Ye|������p)6�X�X|�D�W5hR��;Z9�R�ܵ�	\�ku����[WMq,��1K3EO����W1U�M�$��2-] ����"M��o���dc8j���Jlk�R�X-�#�z�����i=�S�G�[����T|�\͑Z�zh�6�֣f��@㉰�h;�����g1j�LWŽ�.�}����[QF���1�af���J��
��|�z/�*�^#l����>�3��J[ g�b��(�Th;����rIit���.�ҩ-,�v��YI�0O.����!IJ��N��)4�Esi���'���ˌ�s�P���Y<$Ȍ�#��v(�H��4�Y%�RU#�v+lx䃗S�q瀧:7�v4���EV��8Ij|v����]�\³��L�#-Fk��_[����l�7���ћc�o)�֣tSc��RE5E*a����Tf�{6�'ȥ&/�4�&^�6o6H���=9�?��o,oϣ7ˋ���M5ʗ���pr�US���Q�g�4)7�O�ǹd&ȑ��m7i�ז�'�v ��e�y��S�D�����w��$X�R��M9�Yn�]���%�U�
��~Iv��M���[�..G\k"�%v�Yb�H�_�K�˺��.i%ZHfI�C7�	�V9��D�gZ{)�^��x׎�b2nC��sD�'S��mɾ�VYgC�;�Ԇf����O�m�(?�g��G41��B����-.�pO�ڷ�ٶj��-h�щu��.��ѧ�j�o��NMz���I1���J�aC�M̳#�X|��]n����B��>r�q�i�u��C�����:ah�%��S�M5���vg�7__,��c�uT�X��$�!���c�\V-4֡-���ȡc���z���o��wq�T��.�\?��]-��%�Ǆ�s��������T��.�Ҫ���U�	�P�w�"�1Q�e�'���r"\om�(�X��[��%�ș���D�BG���r����`u����-6a�w5Tg����'�m%ύzr���9����(&���z�r�u������[eݕH�EnyMX1����5kɬO_L3౜����*Q�l �ny5�V�h f���d��w��u���uԠ�Ԑ}B���#��V�I�āR9K�liu_�� ��i'�Ytn���α�j����?�*S)�f�%τ�Y���.��-u�XB���I*e���ɋ��M������\*г��Dz���#^$O�	]Y��QZ�q�w�5ӹ��ۼ�Y�׿�We%�q	I�o��Jظ��%���;���Ci�X/�>=ݚ'pEޟ��$�c��9��Q�9RK� 5�ꭜ{{��i:�3������}xRF�K]�0{��襷�I�����č�>K���������~W?<�>���<���������~���/��_�{�|�}���PK   }Q�Ts�7+5J  dK  /   images/6c71542d-16cb-4630-930f-71c4de5e1144.png4�4\�����G%�F���w� zｷ�e�D	QB�����+��=z������]ks������s�Q�*�xؔ� O^NJ��|��` �_Q3?� y)q���m>�Գ�LWm�5��G8�� ��0P�����h(_׎��hx���๓}��2�Y2���e�`e�e���Kw*�/��|b��G��,�\*k���-/X�F��fg��œr�z�cvvJFK�G/�/i�)m�b]��8�X
�LTjYx�*?>��98����O"2����.d+E]r���q��JW���5,�3E�G\w���_����� �Bĺ9���� !A���7�D�L�2`qx�^2b��z�-|�_�Q��o���O���|�w��o2r|u��؁�P,$,��~��v�7�5==�ʕ�����I���1�B'x��G��'�w��*��#N����G�vW�)�S�J�К�V�%�0�=^뽌�S�13�E�j�^Tj�i�xJ,_3��������T��ٞ�Rd#%*1]{<�+KSH�������`)\�}�^�X&.�.C�f"��#Dj@���a!�B��L ����ecŇ�X�\_@買Ox��-�C�����?����dʲ�J�qQ��s�JC�е9���tx,xXb60u	Ȳ�l�Lˢ�:�l
�Ð��ق��}ǿ��Yn�x�t�E^�M��x��-G���M��άG8�jε�:��C��#�,t�H�M�Q~O���Q�)��%#�!���2�cS�!)�����k�l&m��%�� X�)�t�琰X2�_�N��DE��W�������(�]����R��TI��F���Q��A	�
��)�)/L�<�٣�п��yR6��n)R���D'�-�G\
���FF�K�Ă@g0�/"��9�	�M�#'�9H�a�
B�X
w>KF�"	�|s��/iIġA���a>)5�:뿦���[:y"�B"����N���/$5vq!��}�Y$>��X�3�CF1�y��h9�T#���!� h��+����ގ\WggЙ^�E�-����]�ȂrO�Q�����#���:NSA�Q���|Y�,	�����Rj��[�W����vHpc�z/�4g<QZ�v����&�^�Vɭ���a#���(�|�D�<��MQ�KO�Ѝp�/ �l����Ѝ �d+��ྉG�O��Q��{��ڣ��u6\�@B@����0�g���㒒��QF��c��
MHBQO��3�V3�rP�� ����V��J$���fvf�����v�Y{�{~�Ű?�������E>�=d
�=hh����I���Ě��$�/����š�6�:k��D�0�U;��`�e��gV71"�qq���O�,�ظ������;َۖ�E#�3�=乚����ԭ9LZ?�˾nP�6��e=F@$���'�����`B1@���a��C��4	M(���g�1�Kq��t�-_��,����pV��7$��铂��u��)��eɌ����=���m�������II(8=33�Q~�˼F�~�/�g�K�PxPI��y�6n5[���i���X�O����ߑ'���'�à� �����3V �
��F$j�ö}&=�e(!��s��M���&8���(Rjal#Pi�4���O�>%�|�jm��7o�s۶|�-��w�}�7���aގ9��xh�r-�H�L����=<ʪ
@BD�j�C�r޾�5ȱNw�#[�S>Y�b�I��������V��[���|�b�����=_�kX�Á��FpI�����V-��-y��B����D����^L�4-�G*L����pz�1��
U{�^��6)#g_L��B��['�D�Li:�aAU��ɚ�I�I+@����ދ�4��ޑ�-��؎��M��L|A��"�É������ҧ��T���}*�#O֪�x���ٿZYZ�>�$�������~�<lc�w���]��TW�Z^N0�ZZ2�̇ȧ*�p����;Sc***:����hkk��^��?�%T[��;Ș�������k��g2*Q�����I�ʲ�I�H�(�D��mN����7���X�j����M������(���Qn4t��Q�����}���������@�?�̉������;��&�wڷ�����ɰ�I�m$���2*ʠ�:�Zh=�MX���e&���C��X7 �Kz�G���O#����６|���������m/?��l�"�
tIr���$=�е����_��m���C��^Ӷz6��+^���-G ���%�"O���_鱧%��ώ9��r�!����d�; I���|8˗�(���8���EF��׎W{>��Ńl2#֏{��^szdM�FD'1i��	j�V>�*)Y��yq1��8�	��?I�Qz�C$:��h?�􉅲�_vb/�� b?��m	8*�䍳-������@�{��z���ͪdԹ].��;{���X/V��_�*b8OP�(j������̱K�w܌t�Hjz�:�����Ҧ�5�m9���O��Z=,��X��\�����}�W)m�����CKPe�PS"�N��Jq?WgG�v��kt^E�} ̩����$�R�t_2��QRRv���!tZ[G'x�G���| � ����˥֝�ʳ/5���XP��R�/x(&�ݟ� ��xJͣٴ�[?n�|��ܪ������l�bZ���;o(�5tx�b�x3k��I�Q��U��c	GD'���!F"�Є ������}���8��BP����4f9e[w�o��@�l�&��E�1��p�˷�HQA�ֲP��S��P���n�"%R�Q��\ڐ	(��ۘy��3������Ue;�?�u��)�-p1w�s�Dh~�	���:��;J�VF,FR�}�B�.��Z�Q�g�9���O��!Mr5^Х*V�غq�}�g������d~�xA]����H��ː��w�Nf2 c����R��l����m��]���oyےV�:���i5��D9�1@IYy���X{��>ӹ*����D|��w��¾6}k]�5a߾PI>!�(��B�d�jg��/��P�U��\���l�!v-���1�~�{	C�����7�tp��ফ���T�|P��?�DL���QSS��8bBt嶫������~�������*��[�8]�Ă���$���[m'��4�:i��zP�$E�o�/�2&�������Х�'��:E��,�������l��H���g����=�*������3ܹ`J�`�5'���cD�rN�k`��[L�p��& �S�kV�g��� ]��^Xˠ�;�#��G����4;<��ߗ. ���\ 4W�	����2K�n��vd�L.��x�����e1lC�~	vjЦe'A>s�����%��X������	�+�`������S�8q�Ý~�tgc�܎묎�������[��?����OMu`���3�tߑ��v��۷M����}*�3��Z����K��n��9��d1��>6a����\���YZb�Y�閙�%�2��td*���%��p鈈Q/�����R�_j�HQ��%����k�`�Xo'�VͶ�Gn�;:�+kD�<=�̬�`Lj*���&➞~���lUW� ����4��������*�2����m�������vH��"
��UI!e�N�<"ȇوHq�^��UduW+}/	yo�C.A ��ل(AS�
���+���h���J���}�vCF�!ԓ�H�a�ޤ�;����HRS�уC7���rMC��a@F�,��@urzH��Z/�Ns�gK\ۇ˵�.v����/�4 n�pr&&��DP<�<�
�e���5FO���3UТW��U�~�m��� m`*������z�eˣ�g�>�GF�1	w����o���smJ�M��"�?o�u&T��2&�OؘT~_�=�>s�Lo��K)�<��{ӱk�baB ��TC{���o�B@}�ıi���@�FEa��Q V��ؓ��f`�G'&�LMQ�HOO���`���.�é����F͹�F���F)ju_6��4,P�<!A�e�2���m�Ȼq����4e�����%	MM �� �&�Qr�G:�ذژD�K��@G�ϝ�R�u�+@�#�i��b���Kf�f��M��[����=���q.Ȭ��z�y���9tU�d\ò��pi�xAj��-@�'ڟ'f�	������g#m>���J(�P�:��� '�p�bJ��$�9��v���I�(�����ųv�w�^w�77��1�(��Ǉ�������ՋY#r�J^� �����B*cTlB���
����7n����_�?�;oOM�
|8�ո�������BWM'2�bآ�l�C���+Ε���|�����H ؎������X;ݷx�.L���S.@-V{"L��!���+�ao愯i̹(ҋ����F���!T��z���<�l\U��?�� &	����7s�	�'[[[+�(�N���Kآ(9ݣ5n�|�����ݍ�F�o4nXё�̩�JJ�6�pL�I)����-﹠o���ѿ�ҋР�]w���]�oxx���΅b��w�Q��\`��5^�lu;�m�]��nr�������|g#u5���J�|��*7�\^�4	������ Ȳ��_�)��lO$�=�>��3�q$����������9��ZT�Z������^h�?�pV ��uϝc9f�铀IA�#�� �<J"_��"V�L{Է�o��6"t�A'z�#�}}j�Y4�&���,����Ö�Z�rLB�t�;��r�m��� ��4d�����>i ^d�{�}���H��!]E�Y���]�499���x���g�2�����H� t
y�f ������:��Z��3%"
�L�����>i�>�T����������5������I�����������T�Rl�i� �N���W�0 :�jjL [z�&! �Wt<�ӊ��M8�"m$����g}�@�d��N�?�:�	�2��p�~3�=K!�S4?����giee����wfQ޼u�Vi���l�3�Q^'�X�r��PN���F�ÁE՜�z��@h����v\ta�:��RaȐ�V��Ac���*�'��q�l�d���l����2�*�����}���J����(���dA�镑L�F��-u��	OX����,���ud%#�x
��s+b-'�tr7S)�O%V@i��,�3a�;�ĺ�S�����rCRGa�klW���$�5~|wY��o���}}��y8wI���P��e���;��o�,�7K�Z:n��D�UZ�Q�ܾ�|*7��1k ���@z�6 �'I���a�3��ˁ�p�0���56���|��	�G��f|�Ώ�3�;���s��}1*�sZ�䦘����rJ����F%��960|Ռ!�.��� \J�wv	��Gq�=B��ڕ��$i%+��#�����N�dR$
���JJ$��g]�?z����)o�����u�ou(&�u�����t��^(M�:���gֶ#��
dW��Cǃ�b��z&�������l���&i�����dɎ2��MQ��//XT�p�7�2�Ka�Q��4_���hblPmCCC����9e���t7��G ������A���;OЋW���X#ڎi�ǧ�J,��_?�V�<�D|�'�����v�x������/��� ��9����B�Gd��O�C��^���İÓ�k./��M<�8��w��yPp��`.��A;]�������dnY�fk�Z���-�tŭ�߻zX���j0;5;;�ے���vʺ�^��Zߘ�Y�e��b�b[���6���;�u�j||���3pq2h���<7%�Z,����籝����~��R�p��(txyŔ��C�j$j(����Q�t���Na�?�|NM���5_��U*:X��@�c�#7����{	�H5��T��������:i�M�����%{<ʒ\RU�a{�0jj)�,�*�^`�^�b�S�	������W�>�P������n���o�?�;5����G��l_�m�[���2��iii9Jf��])�ÈH{�S|ŵL"^�vtKZ����ﾱ�,?z#��揞�V xŗT�Sm1��r�+E���B��I�E�/�[�����.%���QLw����V��g�{�-�>�k ����=���;��^�cit3Ӽv=:j7�[���q��MVK��Q�I����*ݶU�w ��H�G��4�^K�Y �0�]��8J�z�kɪ)��6j�N�Rl�6�5��y曫Uf׿v�L���x6:4��Q��~������P}����Co��<�6~Jg���ĒF���/�?v����|U(K�����2"bʑ׻���cJ<�0!���fl|�+�I?��\rc��?*Fb��q�i8�iY:������q4ug��c �ɛ��g��PSQ���ճ�j������.1*.:J3���H��.�����%S�[�O��p��i�f�U���l\�������� ��p/p��6tHי�+��!F��9hu����x@G�T��ళw�5�� P(]��0�����6_x��XʞN�\V�:aX��|il��3�<}�ҨOyO�ak(K�`6:l�GZR�G3��(`���'q~�/ϰ,X�����n��Z�m��-�F�Cf'��i	��Q���g�����Z��PYM:������o�
a!���Xt%Ҍ�Y�R|
� � \�����D�_� �8�j�N��jt�迟M(!��S���cn�x��T��Y�V[3�[bƗ��R���^&~~����.���n�.��&���Y��ZM�e�q[�&gb�p_�z���{:��l�K�I�g�x_K�?w���4CÈ9LW�غx]��B-t��ז4�)��g��  T�II�@1sX�?�To���Կ�2���cOլ��$��U�&��e=v�5�K>;7H���~*�j��p᪴,n�o� ���w}:��YD(����J��Ƌu��l�*=�lښ�1q��&"��@B�͋�J�2{A KC w���U9�,9�X�$�����,���!���Ð�ȵ;�]��`O#�$�	\��oJ�	Uy����N��G��.�f�P6�GFy%4=>��_ez������E�m��K�KV�d�MnV������E���Ӎ��
��3�]w�:�g��d�Fv���7�d�+A��OfC�DD�z����ĸ� �`�xj�B��v�����H �O�BAv�zd1J�[�Ĉ�0�]�l�~���3F�0�H1��Ԯ���W{v��d�T�
�V�$#�M,,��d��(����lwƐ�*���Z#��������y�4�rؗg�ۣ~u:�۳�y�m]��2�`�z_��Ȃ��r�ni�����7J�Z�t���}����q���#~�z�:V�ʦ+�����3����
j@�c�t�r�o߾537��� R��'Q�Q��?��dLT
�opJV)rY��t����=�K�;ep4_¢C	rz�\���}e����1=u����V�����x͍�<�0j�:HH�D^�BaHj*�����A�r���7:���߶�$7�g��������=�=Ze�:Sy�j���h�s�(9hΣL�gJ��ͣ�K@��K�i���+���IBUm-0� I�<�Uʟ/�~Y�f���c0+�m}�ݵ��h���r��� �bQ���P�`h����&�72�_�6V�~��J�Z.#L������b!	Ck��?��7���T�Cub��ag���<>����Β�_�ڋ�|j;Q%��Q��lN/q��4S�^��������^ ���Z�^�|�H���䐇����	��@���8�����O�@��\1��_�֏7�q�p{�PH7�'����͍�Y�n�l��LF�����+���3�G6���c���#/�(0[���t���nZՊ.�՞@�Ej�Ɔ9	�5=@� p][+[cY>��B3�]����$!Ќ�h10m�1�T�c�OY�@A}�-1������^{+���|�j	���N��w����Qm��{�M��<��c�w�G�����������yCG��J+1%Xv�L�N�6p�����H�����>j��l��I�2P�_l!�G�zz�9u\��������)�r��`K@֪�+T_�$������#H=H��%C666�����*�ХeP�D	�xW��V�f��� }���ng�Y�Dic�8����� $M�x� ������ɂ�{�?�{�M����t�&'U�c:����JS�q�^�O�,x�#��
���h�������C���%�WX�6���{���s�Y�Θ쌊��:i.�ä������NJ$�HtX����q�*��>�NI�����6VH&1d���PRr�CrT�&��U�?5e��D�~#�|lm_�i݊�Z��x�A4�RU6�L��PLe�=M2Е�6]߀:W%e_5���ȼH�L����V�`+�:h�@�ϙ�vZ8�kk�Gal#��D�������.�?�?���� ��gӟ�����
�t�9��_�%1������9kʐ��ߞ��Bm��B����0P@H2�|�,��i��[�?o/�H���P����:��Th_�E*��H��:Gw��������l�
�fl/�c�����W>��~]�v�ӳ��>ߌ�
{���[q�~l�I�՛p�Շ�k�Bov�JP���4� Bh�;MO����������c�($����{D��������oo>���:�����#�1a��r�����M��G���8��`΁�U~|́�lp��)�q?C�cbf�jm-�r�IR5�����u�ad�1%xU���;���>< ���װ�)x�viG�5�P��ȗ��c�S�q����\�t_�_\���9v�9���$��	�7:��?�,�
ݖɍ;��UJF�Nu�](��-��'7{f�ֈ*�uI���yŤ`�c�/]@d�ԭ��[�h(
�ޖ`��`;�Mz�������xL�>z�ߎЭ0Hh>4��~7�qZ
	F������dx����Bm�ea�j��f�#��)�sU�?諔$u�H���py�b��
�ߧ� H���4R�a7�13$�(s���φ<g�;���Ҝi��@��F�·�'G2�K�Ee�aL�Vԫ��q�� 4���e$��ϴz�s?ap��!�&�ρ{�o%*ɗ�ڭ��qli�? 4�}�*�������[#in�9�D��)���n��li�{{0Zځ��s�֋_z��&�	ӟ�Hݲ�*��F��U���0}'�%%W[�y|��gKf�9G�Ht6P��`��{g�z���&75�8�.�H%e5hn�r�f���f�3i(���E�T�BW��#l����?4^�5��l���B��p��n1H<<����p 4���v�"w#0���4�7{>�1{�j���cs'��I�~��*�F�,m�А�Cԙ��u�Xp�C��
���jʓ����T��6xs�X� g�� О�4����X;oP����u~s���`ݲ����^�Y�c��@�y!���GP^�\rXF��B�+C0Ȝ[�)j�|�q/�ە'�%A o���I�g��Y��VU˴�`�%��%.��0ժl2h��P�R����ro�Qo&n�_+�}������U��G~�,����kzv��ȡL�?Ǡ���7�T�v�N�/�����&��j��p�Y�k/�7{�;�R�T�Y�rA��r�pp�Io:Ͼ2:�w���hm���A�BZͻ��a�Y���^_Ћ<-i��]���s{(س`Jn��P�B��~d�[i�Z��P���˞ж���q1���g�c��*gXQ��X�gϤ�2b� ���8�<B^Zp�iQ���4	N�|�5b�2Ijel�W��P҄����3a�hfP�NL�;��{�n"��f�ΤB-PE��V�ދ
��y�X-Y�l���ڎz�]N�7<���v�n�ta�ڃ�5���M+����&\i^,S� ч��`��C�Op����V�b|��7nXuL_���d���;���������_
�}`#������<OH��0�$�u|��$�Ўc��� <`��h��,�is�5��q�#����?��Gm䊊��F���W:Q�^�:[�`B�J�Vw�f�I�ƛJ̋�<W�ͤ�6e�{����{cƸQ��2��|�G��]����h��síp�DsD���ؾ�nw�՞����NZbؖHZ�v�W7&ڙ;wB˴-Tv�8�m�u���-VL&o�g=�":��+Z�
Y��$Q���cF���`=,�$��:_���(;C��%�6Y��B��%-�k�=z�}���~�%̹F�/6� �Z�d�ɬ\��?)O�����A&>u翃�����~D��>��Aƺu~�����ľ�6��e~���v�qJ�r�L�
҂Q؍�G3��`���ц���iK�|K�����w�����_�-��r�v=4��~Ŕg�1C�\j*�|=ެ���~�aB@�q�:�w�!�p��u�����Z1I�0��|q8T*�y!T�>n"��l���Uѷo.�c=F(�s�-�L�[�x����)L5e*��l"A��j���t�QE��ԑ��,�LQ�Ӆ����풆��w�6pn�_���!#"�.y��i�i���Fe/��,L��)�����Zef�a��M��?��$��.�?�p(p8�ej�=�V�t+��+�f�+ �����"�u�`�yM~�/[{��٢�]�^#��6�{�w����c��0JJ	�������qn��.���@}p�L�AV��O�g��4*�Ǿ*�� )9�G[?S���
c��ޯ1�ӨW&{��Z)�D(gH(1r|�(�^�<�����v*��4��j��i�F���\(����t�5��վj���$#�ԋs���@��&��������ٳ$�`N�%�`.Q
�d�VT������/�*�:��-�vۙ��K�f�X�/Gт���d����	 ��glI���uܯ��t���$�����X���r��,����L�4��u3g�kx���Y���57�{%O���@ӵ�W/&�(~���xv{���5<��PH�ۣ���GWA��C�8Ge�k�\C�̂&��v.��L����r�t�*�9<��3T��L��>{)"r	��$((�V9���~�z�P6�|D��菣��/P�12�Hb��T��s;3
�)�Wy]�G*��ٲz�&V��){^��z��g��t��sI��ή��I��V��-29��HN�6Ûq�(,�A���M��)JJր�Z#�H�9ߜ�}�n�IM��y�wc���[���/mWݯ����I����޴���y�vQqN_(i��Z��Y��]�����ۚ�G�D�\f L?Wv&��ɷ!��浉CEƵlW����/��B�:a\��}��D���|S7��0oO�����������B��7���h����V@�xp�;;�Vnۭ3�,--�	�$��:�ٞ�(�ѣ���~q�@�����~��(7�Ǧ?�T��� L�͎%����&;J�F!+�2%��e���LCs��gf�(�a��t�v�^Vgh�����9�MO�:����Pi£��q�m扖�ǳ�ǡ�����S_7�)��l��&r���"z���͆1��de��'5�2������.k�7~�@~7�t����j+5w�x��ߢ��O�lj��!��:eyڧ�7vN&9�ޛ���R����(`q(����D�M��aTk<uT�@�H��U��N�g'[F{@ª.Y���?��QO�Ƭn��gu��3a��r
Ғz�UVB�@��jo�$�l�����#:q,ܡ��+1IM�T��w��sQ�WY�����"䉖��gϤ���ذ�D@q�)�R��)>x�oK��"7$�tR�g㌽�*9�T�̥�����3�����=Ѣ���%K�__J�Go[ۛ���ѻ����N����;濩��sx��U�q�u����o d�d��֦�گ�M�G}eZiBJ�`v�W�*L�|8��\��⨵�������"==]�|���y������"��V�a��_���<��>~{�z%���]�:��%�����}�R�㝂���G�5�������U˴�v��>}J��s~��q����*����[N8����������G������5�ט�����*��š�����_E6��*S֝��8u~�G���#�3�P�y��p5��Ap�8��?Y���
��������z~�2#�"yE�{S}��2�{K�ǲ�������>U�����C�t�D����-a����Ɍ�-�/_>�=L��X-#�ksg���|T�k;L#�ʶ��`����E+2��tt�DO�����(�o
��a}_~�[M�	]��a~" #(��9�s!lޓN��ܝȲ%η-��a撓g2�@���{A4	JP0��r�d�YTՍ�/�����Wd,�o�v��Vzmc#�
�|�츛]П��:����WÏq�7UTx�K�S��?����S��$�I
��@A��h �\Π�!�����?���t�!�A70j���a�w�� ���=�<5�=ts�%Z�ps�wy����F���Z�N�
�^=?�Ӟ��y��m�����Q�iHA�r�<o�q,���7KsZ7&D`5�#]0չ��X;�_X��>��!�TzЋO#O{���d�{�C<w7�1�{*aK;����
�V2p-GY�s~ε��|�f�5Ϙe���=~���&P�ǜ�?�We6�!,W?/C�T�b]�C�h�%*B����-�O}7(#N�i�։�;=�R�ť��hAƀ�J�8����)���4�J�e;�R>�q��?6��)���ӥU0?���,%���O�e)C�.�fE� 4AD���5%�`0�`�=H��P�4F�jҏW���#<??�g��k��1���n"@3O�\3���TPv�hh�7G�2�.��Y�E�`"W�Ö#�'�װ�I�<� ���#?L��5Y�?r��T���u�җ{{�FPi0O�C4fD���ׯ�֟���2/pE�Zu�	-*'��?�
2�VJ߶3��WDA0�U�K5:����c��\���/>��=�a���P�p�)�o?��Xr8>���"Ab��ƾ�_��k��KɃ����N}��o�lm�o=s�`�,���-����L�Z�`��_���Iy��^z÷|9=f9}���8ս�!���a�Z�E&o�7��T�d�W����I������!+8���u
2��?����< VW�g�)��T	��v�פzm��!@U����o��-/@�+��4by��?%<����r��,��N4��jn������P�����~�oi��OA��{����k�k���g$�6�ms���R�#-�I�UZ��۞��=�Lh�B���m��yO=--�3�9�ޡ�Z�c��v��F�=�Y����K	����KBT�y�Ĭi.	D���0ϖqAǭ�g�2~':R�?���T7-�I��D�g	�	�~����m+�W�"�mmvgA���q�6$�Dr��ZA�lj?fE�<�_.	^���u<������
����z�e�Z@�+�mD��#��!u4��`�⒄L��뷁7���7<�,V&����쾇�[N>����l�~�+�urt���U�{�$t��:�ʒ�%�����ր����Jn��`ϰ�e6��w�~�.��pcm�a(���&�t^�_X�0Q��J2�R,f���+M��a��<b0��6wnp�z!ꈣ$#8�]�S��"���8��R���V��!�\�e;??jѻ㡷��=B��I��g�)L�����lYu�ė�Q����C�/!��ȡ��UHŒ�S�WJe�,����:2|Y�-, ����`����^��̞���c<
,�?
�D���g�^�^���w>��T��Oq�9�A���GK&5�i1����-�)��1���� ?w��� ��O�Yjh�0��#Tbej'�ݡ�'��;�|}�uR�l0����dxӵv,Xeraa9��L_�-V�;��m���jIɛ&w;D�/|��q�0�}����P ���[	�7�"W�F�k�-�7�FyW�ΎA.�Bl��ޚ-9P>����H(<�&spӵ��'�bϖ8s���#O�Ќ��Nq�[��O�hW�V"��]�p�p��N:NBd�5�e8���\t���gS�;ю�i�������Be�\��^����=�
�F?�!�9�ۦ�IھO��x!=����d�����M���k.���/q(l(u�hɊ��:'#a��㫎IOt�M��^|lllX��Y�5����Q:x�I?7�d�&����x�/���ux��U��u���\��҇#���qq8�Ӗ��e���G�k��˥��8'*zR�뇒c��}�/��y{��������&Ϲ;�
��y��.�\"�E��7��Kf�й4����2&+0C/�2~���єPB �H�H3����(g��U�![�c�[��M�d��(Zn��s�®�`��q�.�z�N"��&�v��/#
t�rU+�^K]F�o@b���M$���	Y㬀q�\^�N+���\��S+��_7l��`wWg�)�9�+�\f�I?͢�G�=�t�v�dB$���������\777�6s��>-
" �T�5r��}��m���U�������_O�w�5j�英��*�{��i�q�#t��F����8����Mb�I�Yȧz}��K��ѸNO�@-���j�̓M{+z�҅y�a%��Rd�ɤS"O5��t0Q{>(�d?wy����V�Mi��2�C�Ɋ�������v<��J�w�5,E������`��Sw�IF8<�z����`�(0͇}Χ�sf�ϝ�5V��"F��e���F���J�Σ�UJ�@�� �'�$,���[�����Vx��w�=�9	�[�c���CT~/ũ�1���5�3�0%�P���:J(�w{��&j�"��v�����#�L$0R���u���Ojld.��^�Ε���O��&��TU��z�����'�:ϝ����d�o�|�G%��D bV��*������1SOϴ~N��n�p�������-�,[�Jw�6���a��?֯�ă���ɠHp���+2S�XV<$y������FRD���	s��!�HS�"����Ic��<[��ju_Ҽ�b,�m��l��$�W�gk-��S����p����VT�΅ﳧ��ۣM͓��	׫��<I~�Ӎ�z�������Ht��4;7�Tx�S�Œ��3@��.��i����@a``��������-"Ǐ��$�	XS��S�B�߿,֙�TD����,�xTTT���,߳?���������'@ŧ�|�
g�)ڊ"fn�e>�+U�@����Zt���i�	���
��2�>�Z��,�[c5��~����(/����[�6�kƑ�(��2 �����P�5�{���4�����.�XZp��$�Bb!��&E��y��A�1ɗ����1�s>���y+r=�M����O�c�(�F\�P����5vi)���?W���]:5#�_�������d{��@q�#y��J�N��gg��g�EN[l:M�MF�l��ޠ���g/�l���=3gyJ�П2M��`����1X3��6���d�g~�'�,Z��`D"�O��-��J
�5�3�O-�Y�!~�0%��S*�[��o9��O�9��Z����#OO<u|�S�ɨ^L���P���	d��e��Y'1��������XV���IC�m�\�m$�O���SK�!���=!h����i��;'Ȭ��,�=���A` ]����ܡ�s�+d/fޟ�V8��3T��(Z#A��F2ɕ�}��LP��)���jϾ3y��EA4�ÿ!�I|~��}�rX��V4�=��=1Z�>خ�?|��f�f�.��m������Ӏ@�N�.�M7��xAZH56qJ�e��a��MNid�lw~	u�����`�����T5���л��k�И�������_�6< ��p�)�����N{?\o�p�C����� (�o�ě�)I���Qr?V��d1�)kO�qC�>D򥢽]�:`�^�*Xt\'7�2{4r{I�����_[÷�o�#)�#�Rc��!��sl]�Ti�1��_�҄���P�����)����n�sc�|SU����������ܗ�4�	�t�=��"1���m��)�	���l��Q���F?��Fkw���O��O.��pqN�G[O�gm͔���KҪ���Hvσ����Z�Oϩͧ�p~U��_���{��J�Jq2d��~�6��p��@�*���F7�iQ�`ۭA��8[�� r�#Mg4H��@��XѶ>&��>��(�S�ߣ�!(�ku!|��.��k���?�jQ�(�sE��\�]�ׁH��������c("Z���G�G�:q����C��v�����0'p�3kR�LmQy)�u�&}RU�h��)��;X��;2��� �SQa�p�I��l��x���Ã��k��QMM��k�_嶭���r�J>9@�bs�#����n�8��3�xZ���_�>=�����C��Y@���o�\�Ve�X���w65E���}�g@��� K���^�r�\�ZJC~z�O�� -DϞ5@H��K��D�l��\�zX1���&��CG����ƠT��y�޽����{�{���˘������''���>��f������jW�^E�^��˨V�q���,�l�ZM�y��XZZ���
*�
j���c���ݣ(�ds�ztt4�����7��f7X�B�=��h��]k�eo�M��,K��Ǐ���L�|]��0133�ջZ��̙3سgfff��".��ٳ�/i�F%ۇ9SƵk�2���O��(�3g�qN�N�s�ضoߎ��%,,,�ҥK�w�����T*���֭[�s�N�B�lf����)h�q���4C���ܹ�z��z����E\�x̌������:-�8���(�Y}�"�=�!2ײt���2�og(�� ���Y?~�����_<|��J}��F�W�+�2����f�����>f���oI��i!��9�{���"�ipY���������	���s�d��!8���&�A�)~�3/��h��-�f�N,�P�a^3�܀��̏�N]���o�4�}.K�Y�׳��Տ�U��\��n�u>͠2��777�����>������ݻ�W�7C%$I�Y���H!��I��_��������D�·�p}��#_k�~}&��F^����}������m�=�&02�M/x�e��~ԹW���g~�}�/���o��C��D����+��P*M���{��O���i��1��Z�}���ر����������7�[�g�f�9��zx����^�7�ٸ�|w-�� v�����a����Z�M� 6���޿�9ڊ���1���7l��봙~l��4y_�A��ߑ$�����v��ѭr���)���
?��t���?��?�g�<p������o����A��`@�����GSSS۝��)��3�^��0��g�~1�X,n�i}��$x���c�Q������ǯ������2�ES�ibb��U9�@�ݻ�������(S�����Mp�����H�ػD� &"-"Ph�) �Ҹ J�G2�̬ P��-DQ��0H.����:"��RA=�S։�	@���,B*�[f ���v8�Ի��>�vu�F��o���G��ז1�ވ=  |��NXk�*��
�P�I�:�����6#	H� l"�Oi#%Z燄J 3�Ŧ�[!!2V�b�P��Dƈ� B��rf�B�H$![�u��"Rld)�I����zL*�xJ��k���� ���$Pd{�'�Y$��rb��Ɛ1�����K��r�M��dD�0��T��0�a���lL1SpZ/"!bÜ:�ot:SF�<3�|~�K2ݸ[&+6̅_�7:_��^@m")��(�b���2q��`��Doa@K7�d�D4��N&(0C��@��C)��� h�:M�� TJYf�"�Ř6�z$��Dj���B)Cƒe"%�F: e���5�%	��DZ�\E=P�̖�%
z�w�Ek��~�7zI��0zcPD��zgV�:��ט���F�D�fٲm��S[}|���A׉�E��-=���D��d`ź<�@�!�Y1�LzM�"C"J������Y+L$���T�e�$}�D �DqZj#
 �E� J"���A
�b�2E�$ʊ�$�6&k��E�Jk#�Z�Z��*�tq��Y�~E�;���- DQ�,IL�Y$
�c-u���֚����2i����DDʥ�}"
ED($bf H�a��	��Jqgnn��(������9kmh�i��(��ur B�#;:��8���~%t���8ON�(ȋ�    IEND�B`�PK   }Q�T��4�� ̻ /   images/7a4be1c8-201b-41f2-b584-263fc50cb409.png 5@ʿ�PNG

   IHDR   �  �   �6.u    IDATxԽ	��Yu�yߚ�r�}����EBb��@		a-�ݞp8��ɡ����glI���'&R��l-F��Q�#�-4��@�M�U�յt-�������~羛�*��7�{��������{��U���}�{_�ԩ����l���4��T=�z�z�V6�fsPI픪�ڨ[�������aj8��<�%C�WYH3��L�9SMG�Ri���f�ުժ3�zs��g+��\�R��&T��ڨҪ���L�Q��Ҩ1���a�T*�7G�Q��^�Z���n%U:ص+5��Qg0u+�v��ەJ�=�>Vz�٫T��`���y&�Ľ?$�Rܫ��`��m�'��*�ʨګ�NoП��*un�~��6�Z���I����Q���0<��})�>}Gejj�z�ʕ��kk�pd�[��[��"��ߵi��Zo�H���N��hX�u��hTvW��.*k��h4����a�oڍ���^T���zke0Z�k�cm���T�w�	t7R�V�T봎z�Z�J���H\���{j �:	ԁE�{��F�{��FN^�Zu�- Vp�Tj5~�|���i��e%p��>>T� �c@�C�*�A�WG�����bP���j�_��{iX�`���~j����x��F��VG�iuu��߹\o�n7���Lw�Ύ��̵F��Ơ=Gc�i�����Jsz�`�U����������Dk�����&g�;v�15�ЀKכ�j���T�����!\[3��i¦������;���t��5V�&��B�2=��15�NM���O�����Tu�h�R�sWj��s�zcNn^�sÁ��)8��mro�a�Z�Vk�Üis�e2�'A@7������N�3��6 �z��[�s����V�z���\�]�f��>~�� s�w�)���uoЫ�S�s2�Z���_c��;����*�Fs؀C4F�zc�6��k4�!�i8Z�v��n�Ќ6���:�X;;Zi_|��}�����/��������XJ�45��ިV���6�٬�F�S�6��f���J�V�;J�]0��h��''����si�֬��>M��Z 3��p��� 5"H��J��̠ޘ�WG3��`��]��<U�զ)�F�:l�氚�Z�GM��`��f��U�pjĔQ{�@=ti�~��&U���`ځ+p�8�
��az͙FO�4K�WKM䓪eҲaeU >I�`�4��z�FY������3�Ju�?\�W{��G��M�f��X{��\��{��'kS��a3��ҠI�6���u�oZ|e���C�����-X�l/[�/Oķ��]S������
�.%ޛ{��Φ�\eX�g#6�A�ҨUa��ҥ�+ w������B�A}Dk�fm4���0�y�c�E�* u�l�0�Z���@�� RL�)��-��n]k�괓J�E�W��C*��_�$�V�V�aT�����h!�9�$�6�j��v��?��� w���?E���fZ�p-�!{y�p��L<��1lT���R��9����r�M�
ʫ�`�HC4�Z����v�ta����w�oH���kmG�ѩv���Yo�#�]IW6��a����� ���F��N6��c��7���ԧfG�ֹ���9+)�흭�;k��;����1�r�G0!8%�Ym4�*���pVEXE �OQ�C���R�	����+��lTk��<��p�f��:,X+��&�n��"������4�w��ۂ`�$�x�^��ʆ�+u80����hyv�mD��0����E�H��/#x�� ;�7��K`�J��^!���br�0��Z�F2�]��z�D�a���0�&[�j����Y$}�[g�MB�K��A/���ty����W�6��W*��0:�����t���:HD34�3���>��O=�p�Ȯ�S�.Y�/��o�#oj�Sn���ߓ�t��P�5��O��޵�C�����J�Ԫ�Ȁ�^���ht��F6�:��4C��e�V��kC�^���:��5��� v������C�3Ih&�;̵�-�A����3Pl	�dɽ�l��M�#�qv7���,��[p��F���r��M��i9�v�E�66�m�#��6Z[[c�Є[2r�;v��]$�t8x�	��
��{�n��h<0^x>͂��0��0�?�Dk���]���Ӡ�{���)�huuuH�Ku�4��~���_�W����'N�Ξ9��c��d��h���2X�IYIk��N�CSb��t����T�I/q�#z��Cw��������_��h��[����la_��;�w�{ߑ�f�A��H���F���:���BlTj �-D�d����RZԨ�F��Ezպ�u�0?P
���f�������.�F��0?j9�J����O�q��Y_�N����ⱚ�:[�;x`v�_�V����0a�ܪ�
H���"+�wSkz:-..�;�#=�� �3V�NT��Fء��I�
�l���1ۆ��W���󎷱?z-����\�k&�����M9 �i��4�X�t��yԅ�M'�5-��6A�477�P#%M��fg[�����]�y��{������p�����7�'����y����f^��[�\<�䯮�;��~�k�O�c�*�s�����X�ô���ܫ;�0�:��۽����qe���X߻w����u��ý{�,>�ܩ����Sw���tfgg�Tp nzj�t{��
7��y�|V�m��F7R��NK�.�Y*k߾}���<� ,*�
�E�"�2�-��faa!���H�A���#�͇\T?�	��r3�*�,4�4��߈�m����І��v�꣙���ph�(à�h�C���7a�1�MY5��u�2� И�������joТ��p������?���Ni��S��m����4]z�4��/_�۰\�4ݬ��w��;��~�׹��gy�	}�������������g����y2�DI��C(+ree%
.����ݯ���}��}�.��f��l���F+k��s(#F0��z����~��=l�رX������,њ�� Y]^Z��߮=�cCr�$ph���6�/--%�.)��f�޽�g�}�fc9x�`ZƟ�p�����ܹsq|�����ŋ^���#G���gϦ={�G��#�M_@{� ��`�]����?���E�f2�tg����>�9#��"�W��vف�-!@��>����"�!:�4^�9Q!�� `HtY�Akz�7M��puZ��ܵ{7��;}����Ϳ�7G?�����t����.S�Fp9�y���0=������>���?����_Fpg`������O?�K���-�kQ8���۲���;�����kp�����9x��={`���3���,�އ~���t(/�o�!�v
Q�"v�ڕ�}�8�ٝ�h����r����4����4`��.����>Ŕ�v6�1�n�׿>=�����o��?w�y*���g�`�xꩧ��wޖ��Xg �ћnJ�^8i7����G�&���ao��栃�V�p��=�W���m� "~|�{�d񮝽�ϲ 7{�tן�0� �\��]��s���}x�]w���;���ѣG;$Q=q��G}t������8��8�����z�M�"�����{ϮԚk}������G��ۯ{]j�^��t�/#�S���z����>�K�.^��馣�Kt�s��j�B=�ēi߁}�[^�����鏮v��ӳ��gN������ޥK�y�w>��cvu�#�IX��r-�V��-�/�|��b��EZi�� 2[���r�95d�L�Yw9�~��J�cCAU������`�28d�-h�X�i^�
�uX��KD�cںf�e*�����z��nܦU@�[.7j�5���6��6��_���Rb��VQ�[nI;w�L�N���߾���<�dT��T?�هv��Ϭf��ި�"�ow������;����=����w_�=\�e����8����깳ggn>zs�Knm%�$h� ·��=��p������1MG�j/_�����n��w r��4	f�&��Hʝ�V���݊ ��qX1���8���V��Vhe�^��[��_��&�h��n(�#���� �n���̣q	�*
���U@l:��4��~,���hܥ���_��w�w�툳 �{y.`6-�ҿv��(6#?>��2/���������7�����������y��O|p�"�yl���B�sp��'Ϟ��sϜ�@$x�?/��{�{~�g���O������瞋nފ��������������nk���c��_������ߊl��y��(�Ĳ�#єQm�)Ǫ&���-�ӿ����b|֘�@ׯ��X!V��a#�b��%����q�Ƹ��Tc:����l@��0W�q�N�\��დ���|�|�y������2L���ް�_c^L˸
Xԇ��(&�7�X��U��1�n���GI�<�.�����;��������MGoZZ\����|������;���LM�^����g�=�tgj��~y��?~ꋏ�N���z�*���E����ﺵ�z�O����B�þ�� �2�I��-o~c�5�������^������G�������w=��*Gsp%g�V���YQ>[9�ґ9u/``um��0[cX+ɊП�N�[�Ƨ�>s��9M�nV;�^@\*���?5�9�y�bi��׼��%�l��ccN�9���ӫ䭼�?Ǒ�e(�3fp�p�����w�$`�����(so7�-Ƽxƻ�g�q@k٨��~��tӠ ��n�ߌ �K��K_:zӡ��˗�����k���	��M�O�����ӎ�����G��󒧯�Uү%�K����;>��_��=���5?7;���G?�?�rכ���W:��M;w.<���C����� �D�$��%�
 $���z(\�
�Yc%Hl�c�������5�m<��e89� 7��U��)r�፿?�m��<����<x�������U^�b|�1�Gc��5u�ž�u7��ny��Ԇ�)�Uw�1�����g���x�
x�*�x7�H+i�/��}~�������2��t�w�qە�;���_�B4`�c�~�4?3��U0'�.V>��z�f��Wi�a�޿���������O��ϷZ�dVpQ��,`�B��H���������������������'��1�{��A[fg�g"�Y��B}bრ�����ejx����������4Rqأ�Bԁ��l��)@�Ӛ&�G蜩�aW�}�j/��a(J 0b���~�j�:[R��<��`��/s�?&��++�V��#��X��/�*%��HK�xU]G��vbJ�Yr�_��~I�r�O&�`0���^�
X��,}�6���dI��(t⦇{$jY�P�u��������0ݬ#�n��}�ˏU>����I~���5�=�w�����~�S��,.�D<�2� #Y����Uf�����[<���kR��o�y_��5����?����(Rn�r@'D����_��Ks�|��;j�c�����7�8�,uX	��% ��X)@�+���\yY�&C�K�Wg���CN�����Q��y�n��a�2��N4O.��l2�
@а�g�cI7�<�7w��	�MIO�(�ʥ��;ؔ�IBoq�9ά,q�D���C�L�8K��w����4������7;m>i��Þ���}�L�g�o����0����'�no����='�y��Lw>����.��_{��������g�x�׈&s����?� p?����++��w�������'�����y�Ϳ�ꠍ��_����ן>}��N���X�`��@�E�簞y�=j<�#����Xw���\}Ϡ7�Z����O�{ En�'�{���`���lq.����'ee�a�'�2>z�e�ў���vYB=��3��%�|�`h@ή���IK&P�wpB1&�L�E.�q1���0�d��g��W�/q|�=�q�:�YTV�ɞX;ELEAU�6p�D���]Y�����S����<����Q�2�W�c5��ݲk��?�t����ľ��o����w���'��?�!&2��(���w}W���~`��٨l�}Ӈ��}�)�i3���2�fP�d������.mԖB�_86�G�XN���/;���P�A���I�ͺ��B"��Ńn���%�|�4�������O�K6��Hs|�'@56 �~Ez����t�LZ@�=��n�_y/�"jDb��-��%������r�x��U�7�ǶE�.��ږ��
�29J����n���t�������߶�4�n�	6�c�(�م{�6p�ʕ<pח����}�o���~�\^^Zt)�\/b�^�-ߜ���w��Fgu�������_��ĉ�Qߔ+s�����11�`ʰ���O��$0� ���GN' �2��
+Ŕ����U�ygu���A�+�4�!E�٘��`�|�?b�*k�
�W���d�1y��q�x��J�Y�J������8X�����U�s�tuf�ysU�����w���iM��l^��0���6��w{��T!�Ὂџ������(��͙Ji-7������|��e���Ѵ!��K˨�w�޷�o���+��4�w�����С���ǿ��}(���]�>�D����8ל�;1�X?����/���3�Tv�H�n)ڕf}Z�GFEۅ-,̏�.���b�5�Ӡ����.J��ݻ\_�ɻ"��H���ߊr�������&k6�Xz�ہ^,��Y7A�����+�Ҏ���ɘu��t���� �"]� ���}.��v�V�˽���b��b�����/å�����"�嵮�&{e񩩼āY��Gx�Ȼ��{.���o;y��#��Ǫ;�8���Ղ�-_<�w���kZ}]�޿��ٛ����g�y���wJ��Ξ;����w������w��?��oy��O5����d�R� KL��<���h��I|�R3��$Ga��G�E���s��n
�r%d`h�J�M�E�֗�5�|en9���qF�!���6�h\d2dp"@� {^��bS7�'�#�JT�{�I"���1�`����C\���O�1���s�{���|�� ���/�mҮ�+~7A�q�W�"��|��޽"<ޭO�C�}|V�)�ehEty���w�yw����ؘ�����g^���zh^�"��lk��YY�y�7_�׾���������F�y�OY�������Cϝ~�飿��qЁ�3R��<�����Rg=D��st��e[����	B%v���<������>�G(�"j����e���d������g7���䃻`�ar#��E~4���@w��2��JQ� d<g0�-�ρ�/��ǱN��8�چln��R���pԜFx��4�^�I��\�&�9�����HW�޻i��՟���=�����{ｕ���ﺀ]����Y�� tn6�'�X\h!|𶩩�S++�U�k�d�k��>-���ɓ3-�E��D�������z��������/}�ᣮah�X���y��Ƅ��
5�ᓐ�� ��V��4VeT1a�G�t;rǜ?���9����@��(���������E�aۭk���b�Կ~l�=��v"g&M8u����4/��bW�ѳ�+�l�ٕ���:rJ��\6�|݆[��tH�+N�����Xp��"���r/f�k����t�_���!(�e/H�ۻ9��eC׉u�]�|W㰔������ df��=����Աc���_S�?u0�8�o>x��W5��D7l���<��{�a�"9�v�J�����0\9��c���W��ڣ���k7�v�.����]2����\h3�ef�AD�W�#L��o��]��sy7�b���m��e�X��\�l3��Ï���h��ޏ�j��6��d͉�[�R�\b��a�n��Xg��Bf2Y3M�`�x�����^N����`Jy�t<G[ۇ�m?湔���Ky6��>dx�    IDAT����O�O�9�g{݋�ڌ×1j���R̱�l��+^�џ�ٟ�\��$�&�1ק����=w���똼��:�����W�ugs�{#�i���TR�Jܷwwj�����4`E��e�Q�VY�In`u0qiy)Ů�̳6�-�6�☉'A� �LC3I��.�6���~��C�IT�n�aC<b����iw�x}~��cr.{1�bm:|���74h<�Įw�ʺ���/������n#f�����8^8.��z�N�Ӣ��nᪧ��t�t+�%��I�W���,�Q�z/����d���nw�L��/]��L�!q�s�������_��_�x��_�rՠ3���?v�-�^�to&��'�����2�|m{�����-Dk�klXJ�����+��8nip�����T� /�AN/Q���bO��s+���*��ƈ�5��P9�w��9̤=��dw�KT/�-�4�	�{����i�VByqe���p�W�yg��W��{Y�Ȋ76$�̬�(*o
Q%��Μ��7�]YM��N�>�����p:��P��v����ŝ�m�̯9t֞V~_�g�,��4�[�b���~��~f�~|.�x��~�]���2:{��`���`��UR�w���f��;�>y�q������c�f��?���7��9��G�E�<7�����'��X�����o��'�!���*k�i �6��c3QM ����	�D��A|OЍ�F�FL��_؃�,=!/�z��	b0�?f���d��U��\N�;���r�V��_H?��ߛ~�'�}oL��c���z���;̬�7�k�c-Hħƀ�=������ ڣ������}��!�O1x2=�!��ɁhЇ2+��eؽ��$�^�[�z�Aclo����x��ڞ����a}��ƫ�gY]Ӯ��/}	���i�'�|<T�kk����;23?�.����<\����]o֏*7�(�����G�{�P�͝;{nJ���-��#[��V�пkC�ɀ�Z�����G� ��8஀1TS������?�j"B�����B�i)\<89y��D�=s�R�;?�w�;�y���׼P#J�Y�ȅĤ{lx޽�^0s�e�+�9�!�� ����g��w����w��~��>Ė�+�j6����l��W��(�n�4/��!�F�I��<��:�=���%�k�Z��-'Wl{�G�?���c?�c��[oM��ǂ���vгէ�կf���3�v^Y]�ET����l����uZ��ڕ��Ȓ"c��F�u��r@��a(Q�~՝�0�;�t�W�� 0:jE���c<2���8gH#��Dp�<K���A8�$�O����Jٻkw�����t{#�G~$���X^�H+4R1M�⍃C�:K	f)o�%Ͻ�3"�u��"����^��q���tӾ�閃G�/$;�u�?'��^B�xH(�$G�Ř�k�'���k�y1�M�1��{2~�帓F;/M���cq/~��]	�B`��Jw��#I���ߟ~�~ ����+1�T{��T����g������6�iHC��NW�?ɔg3r<Qj��խ��͹ʩv?�yӖ��% h�W#s�1]"��ݳ����,U��W�^���{L�D0DD�=B7q}6G�ʂ{�?�?�~��~*zOv�ݧ�v +�LM�R��@����Js	��"�2�6lv�Μ���"+�s�3gӷ����w���c���
�|N�=݆��5.e�T���z��I0Y�k�O{��)�-���Hw2|<�G�>���/�|�L��Qc&�����Z�݀����/~1@���iP�_`�Zm���5��=!ou&� �W�;v�sG����÷m�3���򣜫�&EZlp��^F+�xg3� ���\B����! �HA��n��wWgi���Nd�96�J%�F,s%=t�6��\�cu"�I?��ޟ~��ޛ��?�����/_f��q�+�zZ\��a���B�O�G�xfc3皱�� 8�"��9!:��Q�NU@�8~2���#���ߖV�	.^^IQ�'ϞN�◝bI�;z�Ln��c�y/d<���=�ԡ�6(��*NbB�����qz"bO�����u`Ᾱ���tB\���w"cP�d��;�U�+��w>Bw�"ꓞ�Cb6����=�G�%�%r�jS��^P|� u���<�ݿ'�20�ڷ� ���$�z���` ��\S���[V���o�;j����ڿH���:�I�R�ܙ]��}+�פ���yw��Jq$.�U;�ڈ
;w��xn֚�s�A�_~�{g��U�6�)I�R�ڳsGZ�t�6��e�2���X��(��UQ������:*�U� �� ��,�an�R�f{˂�m�4���������|:�z�5&�R����r[Ȣrw��L�������	Ĵ%Mt���k�->mi5IG���V�H�Bs�͠��`�r��d\���	46ƥ1L�d4e�=�=��=�Ju�s��&���m�~���PGG���y�Ec��f�v�S
�I 춞3���eoȫM�G�$V�&��zZW��9U�l'�G��V��8 �ҕ����X����t�]w�!.'\z���1���HZ,ɽ�]��}�|ZcAm�6;]��dznW�8B}�͙M1E��M
�9T;fgL���F+����3�G�T������ԌϞ9�����Jg�.�U�p��.���E��Z��^��T��aB=WU҈H6���Y�A�U����M�n�=ד�'S(�W0@j�$�����'�o���GJ�(Ø�n�5|��a}�4iykLt��aG���I�Q�jm�ڵn�y���w��<qb�I�>0�=��9s�|�BX�R��,h,dl�3���E��eL��;�
�L����g�� -&�bU'�._:����7�����I���� �9��tGD�H���u���@�����_XS/�����`F$k�����W�퍛I��`�TnL�s�q�Ip�*�g��K�2х�2��uy��w��">�ܩ�O2=�����w�5�K��w�#��W8����$"4�<�cj!��wa�a��H�B��,�|�n��:-�wK_��R�M����\��/�3�-v�UZ�=D4p�h�Vf.���Vޑ����y���>��K�R~������!���tkz�aW��Pg����=��gb���(�<o~b0�����j�R�%�<��X���D*B���kz�h���5�񹲲�J����p�}1Y�L��ƨ�Ђ �yuWN�J��Ҁ��2;��h:jk�����BL�BC�1�x=��"��R�yP�i�Gn�����?�D:�[ED��Ag���e1�-1�D$ٍ۱W�*��N�G���O=\���Sy�M�u�政PQJ�lț��!�Rli�I �n�+\�pk���1Lwm=:�)��T� ;��~�?��������Z�-�:�;��z�'�2C�G�՞��*`ɉ^����MfGjC���AFs3��啥E�I�:��p�(�8�n��c��[�i1�.s��	���Y�m���]{�&�𨁟�'�8�y���3'�4@�Xe��3�	Q{p�S� ���p���rڀc;Pu�X���Ȼ튬��iT�jGPq�/�_�#}B���A��H��M��80���{<A�u ,�bn@���6��t+{뷥{�}]�(�?{�f7���W�*���X׫�0��b�i|[�վ�Rҭ�W�:��\W����D�J�"�M������K��p�˭����^6��uc����/|�~���[���Y{��z�F7?����}3d�A
Q��N��~&���	Q�0�K\>oAo\�lY���� ���� p���q;vK����u>~6��}�8_h�S�{��kp͓�}9�/�O�����Ѭ4��S,5��0�߿l����"�Q��C�'r���54B�;������!_ I����J#08�>��	����[̊�h;쭧=��|���6�z�p�̗K�?��\&����'�oV֖kKK7c��xs&cis�r��������f��>�V��h�]x��lH9��0d4�g������jL1R�J.$sבu��n���+`s��a�x��~��ʕ��F|pe����& �#�k��HX�( Vރh�W��W�L�+��ь镟����M˖�@<+����-oyK�G?���Y��h0BW>�\�s/q~�n&d�?�h���Ӊ�T'�,��ڼ�m�В�9�ީq�lҩ���
RW�y<G��$.E�S��&NդV��ĭ1S�R����O�?�h|���f9.Ã��hI8c�m�i7~j����sHP4I�u40�� �T��Jm�"����(�zy7/ l�.�:�9�W4�q�e+�\���S��ǖ�]{����)y�.>���������ǉ�����upnN���8g���ݜ�\�6��w٧�n�L[����֮�*;�LI{Av�w"�,��rU��6n������/��ϥ{�]/,q$�M)k<��G�F����s���=��� j����i��5w9��	`��\UY�� 22 gZ+��(|X&]D>_ر��E�@�Z�/rT������6��a�3����~�i�H�k⦶D �)�f}*��*��`2�f6�~������v� �RS�C�y�x�\C�vG#}��u��*���>y�Y���2)�j|πͽ�n��g�Xb❚��d!DF���j���l���zm��޽/����p89����B4S��� �%[���}�p�K*-��׮�+�˰7/�{m7�I�����ݖ��?��t�+_��,���C$oʦ;��,8O<�x:�g��9 �gQ���"(׈���@jED��8���LZ�f)�x�7'��a�e_h@�sH�N���K����N���,	�R>������"+�X�AW^������&J����Pi��/|�ߗd"��R��_��y�nU�t� o�{a�����T"_姸��r��^6�F�g��Y�g����n�\e��:S���1���Tk��Ũ�77̹I4F>N�68T�c����f�hip�b��d��f�6	q�FX���X�r	�sӄ�$����3Ǖ��>7�/?��;����'�����4`���g>��t��ϥ#�ȧ \zp� �8]8��r�=��gʕ��I''@�4S�3i�!�Ѐ�j3<yG�H���x�w��~=f�؁���j��`�\@eAN���~6q-M�M��V���6�r���}u,�������S'��+i`K�]���+!��%<����h�lD�VSh�s�؇�Q,�N�r{����f���
'��	����c6s�����ZҎ7A�r�oݪ��O��i�I��������	�L�=E�F͹p���%�����N`1&�x/�;
[(6�/a����7���W[;���E���ۿN����L�?���S��B.?��G����t�-��>��5��2��2mL% ��Tī�Ь�����9����W���'Ʋv��!��@`��9dcW����s|�δ�N#
]^B� �X�iL��-∹�>@����w���ѵ/�:s�1��-]F��F�~�s�Y/=|�Lڳ{1-!�HJ���1����y��VM�4�7	�C�E�V$�ա��2�<gcrح:,75'��lk�,�|�Dw��k���-Y���͎z����ʿ���d�hV���lo���+�-�o�/��F�c. �Lɸ">?V��3C�iL�#�m@?��M?�C�M�;L��Չ����i�w�s�O����i��*�r����. c�%��D�wbG�yԡ�"�X.��+1o ��/���j���������i���YH�j4�MT���Sس��R�B1��Qp�<1p��Qıspp�z	�3�����T��5*D,�^f�ٻ��c�_����Ef3�\[?g�P�c�1�1C�\��ľ��۲��M�1L~.�.I4�N��l��ڵ1E<5�ůq��G����{`�C؞�tN+���$εK1��K� ��(���k��ߟE\q��#�b6[,��b_�`���Z��7i��~�p�U\z�ь���Mm�N�;HSgܡ�����N����ʙ3�>=Bg�d̀uʳ�q�i	hMɓ���zS�U�,����q�v��k��^͛�tz����QE>�.�.l��ľ�H3`Q�"��*.�Jaa�M��ʙ�
Ո��t�|�5�m��ťt������ߙ�Yܛ�<r�5�q/4Y�I�����?�5��+3�l������L��Y23a�~\�>��\dKT�M#���ڨ����67Ĺ�҉v8� �����n���Y->��(��>s��-Ԥ)n4>�4�� ����0�%���~>�t�p���^���Tn����G�U{?Y���-��3[F��"('W�l?��ט�9���rN���s�1p�B�p��` �<i95�;��B�^j�A����q���!�Uq(��^e]>��i��KT��� Xڅ�S�|��o8v';�6��J��%�|��T6�7��,�VM��\�d�����~� >ק���a\�<WX�Ӵħ�/��m���eE�YcsL�5���������?7���m�Enؽ�~5��8�&" ��J��M.�*2lzɅ��AhʩT�7���F�NNeoFăa�f�n�@�'���P�~:��fn{晧ө��J�3s���I��#���Zѥ"��GT�@�2�������L�Ϧ�Y�vd�M
G^qs�߽��*��U�ˈY�d b�3�ӽŠ�M�tÔ8�y�&\U]e���j�(0vP8B���&~^�� ���ͺL���W��N���/=��	��ӈ6�g{/�Z�����b��t/��=ב�����rz�����l�+zD���
Ӳ�S�]���W���b��;�!c�{>�__k�EEO/W�\U\2kf�e>A8V���2��(ﮃƖ��N����*L�G��7����w����ҿ���v��B��b" �Z����@����'���� ��}�tϤ���d��3rx�o�L�z��f߽L�����=%ki�u�s�u������v���3�P��5�c5~�͌'J�@���%�p)�K>�<b���P�9�P��O���#�D,�4n��Aj��F���M�N ;s<�lV�[�I�?��t.�L�-�l��w�˜��ft�0�
=H��g��!����uFP��ɍ���a�Ϟ%4Y�ųV��?��`Q�GYۺ6�b���qbt"�"T(�.̥%���Oͽi	w���`���;���N��i���S�=Ϻ�`,Pf��:O>�>	t߷9��'*����W/z����7|����A'gg�d3L�4���~�QA~�T5��hE�Z�l�K�fĢ����@� NTI�/F\\:#W�n#[��3��ʠ�"{�wltJ���U���Ï�8�3����U�i
=:/َE�tZ�U ����
����N�O���34�@q�=ߔ�L�����ʈ�#l�� {'��C�S��̩��t6O�6��y�V������.PK�J��ٲ˸���|���.N��=}�u�d��"�<C8��Z��&s-��[\Yq�w�x0{�6<�Z�@�]�f�f��]Fk��
��	]�m�]n�z��1�,w������OR9p*����,�b� o0�|���=�;p�.�dЦ!8�)Q��)6 L���C�|>b�h*��;�B7:�1cRn�������\��o�����E>S:m5/gS��
m��(�zQ��I״����u�������\���KM��Px�
ǐ��S�<�q�ƫ���
�����q��C��;��bV���4v{F��R��5X�jg=�+���."����L��r�}�X�\e���n��]cʸK�]$5@��š��jYu7Y���R�R�r/��%�f�m�>�+W ���=�r���MG�
��	4'J�\��~ .@ѿkܨ�    IDAT���i/����f��mqn	SM'0<Mν0�p��#��=ߛ���J���Ui{Ӳ���XcA7�E��Efo3�ƅ�U�+����_ ~�����ao�r~�rN��ڕI�2@��8��q��q]9]YhTl,�o~�I)z�3�E_d���wߓ承Όh����d<�-딾�6���178���D4r�|�-��U���<b	{�5�nK�N��l޽̓v�b����5+��^�ܨX�]-��a�[e�-	�ƭ��~/*���[�R���{)p���_q+���XKN����^�'���o���1��0�OV>��͌��O=�N��ob���$)���h&_������U�jw��n��hɩ����+�Nm@���3�ɘ��)�A��6VH��^f�+õ]�!'W���$�w�1�֘K#���2�&�!wg.�o�3po��Y�z��'�����xi~��4˦��L�_�1`><��^{���矤�6~~�K���.�BN�L˘��xъ�d� �ԅ��f��8���+������ɺ7��.ǖSkWw�;��6���Ԗ��D��~C��ر���#id#�6�9Y{N�'��{K&M�dz �1�^�5ig/My.�aIr��؁\iW�!�����RbwP��S&����g�MSI~�#��QA��=!��q�������m�#P$N�Lm(������Sl�=�� ���Ɣ;u� �ˠ���U��C�W~ﱟ��������ܝ�e�<�P�-]A Y���"��&�ɷP+���;M!&bG���=�qc?P��2a48^x�D�P�o���txa=jG��a�̆�T���sQ��2`�N�q��y���K�}�2��W��O^�_	��������ۚ��wم������8�?�����(�ҋ�=7_f����R��B������l���}�oy�C��v}���l���O���#S.�f�?�m�e���4�� �%����If�����ʼ��Mk~G�^D�/�ٟ��>�.��\�*�ԔAϔj�n�@�*�#E��T�2wpb9�y֓�+8�j�dE�X.�xY�(�BKa�pC���Zk%��(�Lr:ζ�]�p�=;XW���f�:y���M	���8h\j8�7i/�=f�x�fo��8�sWUɻ&��{�����.#�\۸��4�����)�L��h�֎��Zn�!p�l�'S7
�Ի��:�9v��NrҘQ��/�.s�ܽ��hW�OƱ��mGV�'4�wя��w�}�S]�+ru��C=�?��8B͡�jЭ:(� �xT�~��$�3�. ���qR��1f8�!ו��d4ʣlh�T��+L�;Hko��i8#���j��ĲE%�3�̣?�%� �q�+ ��0į�t��v���� O�K\} ����9�P�^��Vqe'�ܱ�{�|��dH˝E�d҃6���U�d}�z�S�c�N�{�a�W]w�uJ\%�r�wq3�Ԟj��y���/�����ùy����t�����z��*�n�*א�Z�Gf�D�ϚRHߣ°�^�����8TMł|
mcz���S�����T
bXy:��3ibՐU��7���չ��9�6N�i�Z���No�����t��'B���n����y�yF�����}w��	�yf��W�bBrC��(�o6\Z�'�hq����co�p��+󦆈(�D6 O��!�=#���{���m>�t�Y��(���i�<�� NZ�,���A�;�O���[��R��;9n��Wȡv�G�bL��u��8}�2{_�TH�D@�t�*��ue�Pyө�h�X����(N�8����yAQ)LT~T[k�*�gk���q2��O���3������[n��@�XR�Î2�X
y�O?�R.@8��E�-��AbG��C���x���)v��%���W�F�md� ���K�|�
p�B8��8�3i�r��q�J�ҋ���#�4��Q����[����Z�ӈ�x����Mhd��?����+���0�<ɦ�U����(�)���:$��ȏ�Q����u�яW�� ���=�O�(G��+J\���ɸ��H�qVj=�zis]�
~��۴V�YJ�ϨߺbH9>���_MJAlW7���3��~�Ζ�&�.ݾǃjv�)`�~�Lz�G�h�w坲���A��KP� we���ݜvt�7����<��vz򋏲����&q�%�6��sPF�!V�8v��3셸���+��	d��gG��R�B�ɻ���+U��
�bo|qR-���v�� ::ɶ� �Nt��=�$���%ݼ�u�g�2~�C�׏��&M	/(5Qd�1mC�~z%���{�k#�VIbh��p��:f+��x��f�Ih�A8�'�9
2x����������)v����ɰ�LBU��_f�ȑ���E'\ �����I�����,ge1]n�*�Q@T �qHe�D�ͺNd��G�Y��H5MsN�i��C���ś��k�J(rDu�+;Fz�l/�&x�[���?�w��4��,4 E����e{�6M���8{�	T�zu�*�m�r�+jq����|������E�j�L"�@�ٴK}�Qy�*�͌l=�>�g����WBL��^Ϯ����r�R�L�,%�W�o܂
}>E^�.7`?���[\!BI�d�B�����ݏv��a���h��]������7��8�	9��+������	&Ťj75%�H���{A�I�@���7Ϡ]`�b�"�hQņ6�M�R�Fg���@�b�������`	-X�["M$8�)�[`Ƞ7�2��F%�n�c�θQ����A"�� �Ac�}��ZCd��|���сY^��!�A�n� ��]7�� ���36Je�h6����z+�.T
wk_��ʢO��('i��1�s(�)>Ðf]�y=s��~�=;��9	1��X�&�٬�<f�
��@)�ϥ �7�cEL\ž�_�o�n�������@A���'O�8-�t��2�3s�>�E�4M]�i���Y���M�z��SMO>�t�Ϟ>�P�f"��RY���x���&rӍro1��\�F'MN;7� ֍�5ʝ��"Ϥ3�ڦ'���lM�ȹ�(u$��l��=��g��L�jLu�'�vլ��x���I�����{ɧ�r?��8���S�;�u2J���<�q]�7��b�t���H�'�+�fƶ�k&	2��]��-�𺖮��4ۤ�=����Τ�#�xq�;֕o��x�=�-�w����dAg��\�[�qڻ_��G�\.�'=���9��p`��,����w��`����+�W�.Wu@�ϨP<x�X�b��B?�!BO�#��QN�J����G?��~MŸE�Cq��&��D�2��L�g.��g�2׭��ix��q��ٸ�Ճy�e�b&ӑQ���ʻ���&o�,��4��-�]�����s�K&<��%�.I���xŋ�����B���|-w��3y�21z�Ç�~���1 ���c��r3Ƶ_8��L�Å��L�Z`X�r)�LS������t��[�Y��i�W��C�"F�(s �J�y0�B�(�؟v��i��'hS�Z�O2������[���mc�!D1�SS|q�w?N�#Q����3��iq	h/M��~J����h���̻v���8�S���W~j�u��y�Q��_�l��K�����{��vB��$K���Ff\BJ��Ѭ�v����K��5o����X�IfA�0��|��f����"m�n�Ҡ��[�J���p�&�$�Y7=��
ʪ��q�XQA�l��G^%)��>�-v쬥�_z(�X��]:��z�xUM�渂4�p!�#�嬔��6Ċ�A�jZ�4Uo�Y�O�sY6�:rw��=hå!����ʹ����@��>c׃��6�lE��{���:*�
c�a�^�	�9D��ǭ��_�Xb��K��]��3��Lk�x��@{JFLs��}��ֱ�ԛϹ�sc-X�R�/�R��N�?�u+N<��g�&r<�vֹ�mϼlK^�����N�WBc�w�62j�hJ�-���\���G~���}ҭ<O��l�eiL��FQ��4kN8/�]��1�c#�1�/?O��t���i��<j\�R�h2�v'+ *�4K�@U�+ؼ������!�G��4J��g�n�z�q��R��U��v�<>?���+V���9�Uęqן4*�+qz/v�^�,�O�'�M>?��G��%.�Q�CQ�Q��/�3�/�z�t�}�;uO9�6�ġ<%�ϓD(�*�(�X���(�fl���e}�\�V�����g%�� ��p6.�C�W���
�\H{�:6���MԂb���v���"�U�g��B
7�3����@�d�GZH !y����R�Є8�2���3%�!�O�9->��`�N��<�Xā��YW����yv�	�0׵�W)W�Ǧ=R�Z�-��{�W�y/n>;�_�.�O���ne$rx&�#/�!=��I#J�fs��4�Z�&:mz�8*p�E=��@�%��^�}�c������]����ɾ��5����D�I, ��#8 T�[��\2�C��U#P �Z�k/ZR40eU��h��2ĄqE(�X���E<%�F_��x�x�L�d�Ы���d�S��]���n�vW�C��(��9zzo��~Eg�����2n����~�5�=�~J~���v֭��g�d�ʵ��Թ�'*m2��g9��lj��Y�s�(5�?���E��yL�YcQS
��@P��F,�o�9��x�	�C9�D`XeȲVqAbL�.�<P���]�'D��j���,� ��͑����R]d
~N�8qt�o�T�m��z�9�oEY���%��(�"å⧔�<���W�6�I��T���\�Phf�qEx~�mO�/h.s	�t�Q�{��'Aܹ��Uc�d��uoyʏƭ[��0���I�4��F����e�kv�<����S�7�ڼRn,C��	�~KW:�S{dC(��t"%�T��&ʜ�qb_�Ѹ�LF�+���h�o� �#2f����rq3���+��	ϓ�RI�ʗn�s;Si�jI���q��(�nu�+��X"1'�c�]��EOd��7��A��`l��Y������]��w��E��2/�[�?y��ڦ�ơ�v��1"�q�tӽ�*<��n"N�1;E-�{�߲K75.�r�jQ?����f6B\RtAl1я�c4a��U)��%���տQV%\�7o�\��f�����c3�R�=3��Ʋ��2fHp���)�'��䙕XfH���R���R
:i��/�p�$������6�-Q)V�1&�D�'��g��j>W��K��	���p\p�yw٨������o�ek�vW�ɉ��+���p�r9�x4K^�Lp+�N��`΍"�&�"�d�uW����ރ��1��z�HO����!��qk�	c�^I�k�盎Jw�~�xL�'�[��l���0�r/>�~��-��>J|宨��l����E�my�#g�q,_B���͡�zy&q.^�Wa���5qN��۵#y2�y(��n�BD�����$����s&^8dhS�Icr_-����0���?z0*P��&�<��6tYk|�����qؕ:�r��KC�S֨�膛���>��<ΨQI�B��ڱ��S��l �4��%F���b�Ʃl,��g��J�n����2ZO���h,�߸������r��.u�����LXIE�F�S�(�n�n���a&�e:y|�{ae��Ϙ����ɸ8�v�<;׵��Fݵ|\���1�v�og�x�-�x�s҄;)�ٳ'�c�� pe��1�Uc��Ӕ�o'�����f� ���`[��J	VTLTkT�r���k˱8^l�{�c\�]N��ӓé9�r�J�AZY��G��e�h��Rc�wcn�*����Ԃ9-t�Ư~z@���v���;�?Շ�P������B�E�z�7�(��vY6��Ǹ��W�uP��H�OmH��6Fp��H����#=�W�����L3�DC�ԏ��|E��3	҉�!��`����ə�তY֠h��ˈL�׆ g�i��ш�ǽ������2"ש_0s��
�\��K�� aͤ�)�;���`���@.v�U����Le�sL���@	剪����̠����$;P�Ո�Y�sx|� ���\�P�� p�X"J�h������i������8g���y��L�7���J�of)0DY�Cɿ�&i1pl K�B�w�!�(�b�8C�i��pDilҧ����|����>f68�\��p�ݒw��c�����9iv��RZa��	m<���G��,�-
P���^;�K1�/X'�v%���Y{3i7N�d\bi��h4�hM���ű��:�x &m��+�p{�neuu%�bJ>����	��Fؖ��Z/��LU?�g�}\�ؗ����m�!�nN�>w߁�|��I
�u��:��YGD`됭R4��д�]���SE��w��;�O�[P�p��nK~��}��1΄N����qܑ��,��	=6b�x��g!���UQ��'	�f̥3��⢖���\���a�aXXa\�H]�A��p^փGħ_�/�(�s�l�L^A���.^����RA;Mq�~�X3!�ذc�!�)X��?�ȱ�<F�+�̤�g���p���V�/�$� K���终%C�s賶#87*�ؕI3 '�[]O������I0�]�+[���C������G�����x���_F"�
� �0c�����G���Blh;��-� qҳ���=�����5�N��'��ES�`ײ�c�{�A^�:=�B|\�5�S�0���p�&��|:\�v!�s�3����)��p6erS�1�H� ġ��nQf�!)�`l��z��(�,�xx|��S�߯/(R�µ�XS6�n!������A����+~J��x,"�'��/��ӂ#���}��K�G}.G�H�գ}87;�)�{ �
rni��`8����%��g�-��z��3L�|���a��sQ�\�xMO�H��̉�-��^����'3���p�9 %7�3�pSzF��4z�~�<�A�nPX9u&��.��l`��j�@ˣx�g��вxn���ß"_�>*�Ԇ��C|�Sк����Qoƣ(1C|��u�)�'����7@������Lm��1��8��J��K�r�i`jn6�O&$Ի�i+�L@�,n�v��i:�& �d�{�cm��x˞����e?9�����g�A�Ϻ�@BQ3 �/������p�h��c�w������")��绗 ���,8�-
o׶�X`�)���Y��׏�������A0h2��!���Y�	��� ۅG~�`�])}�y�*f�#4���8��1d� .#j���\�p� Gu#&8yU#�D�i��DB�H��� �
j9���*���y,��	�d��%�=ӌؑ@��ir��5�=K4�.�q�����c��F�#����{D��+E��ORc����3��o�K}�z`��`�4��LS�h�[��؟��s�My@Qư��g�[i�c��٨���e���$uɚ�{8jJ����%z�Bܒ�R3�cEX +�g)�	'󿆑c�0� sx�k)g�S��$՛o:���
�?�#~����Ө�:��z���tQ��N�ʋ�o�y�ݐ{Q�O%|(��c��` �,�5N�m*�S�~y,����3��Ď�U������~�2��թ}t�Iy�U��#��q�3;�1c��^�g� rA?����� ��0?��'B��':&�G�6kh�t�0��]f���$�H>����q���"�[v���u�U=��&�e����˰d�A;�牯>�2�vݥ%����"��}Sv�t_�OM�%�L���'K�5��w+�L^�X�r��ͻ��n~\���J�RQEbԘ�ڷo_�}���@�.��AX������d��;wO�m��]�\C$�4�s���'RJ�,�*-���=~+�ˏ>��'��)�Ӟ�F�6by	}8eS5����9�(�    IDATw�3=�g��&�Hs���<��_����3ir
GV���7N��UN/ӿ�C��(��ʹK^J����[�_{�7�����n	v
�W�c�m�9�_�hO3�6jN���#2!�q	�`��+b�@.��O"L3o[�B�)���R�Cę������#�.���^@>t�P�g��X���ඞ�z�Uw���>�X���'��/��Q�H�/��a0�"�n�A�z�mX~?�md����yn�K�e�93{����_��:�uv��=�:gyZpw����؞ECq�˜'q�)����g{����ۡ	�Z�GS��:�I:ƹ�p��F'�e���i�o�_|��#t�-NЪRF�J*i�g������J�/�I/��-��ͷ�~,���y0B ��C޶��+�(^Z�>��Y�ʍԼZ��ze���jYT��$��4�����9
O�̈P�s�Y�sC�~��^�P��ٻ�@����Tf!l��R6��@�ZF�P��R��w�h��IS8�r���zF࣏>�n~ű���*i��c-Lϡ��0Ts{w�[o�5�<�t�G�n�A��g��t��G:��G�t�a$�XDðB��k '8��j9 7�7ה�ʳ�=�S���F��i�:�*c�4͢,�Că��Q�Vz�b� �F�=��ic�*^cORz�V=U���t����;�ǂ$ft9��A����Ȅ�~�a�'�H$) �?�j����r��ز͜����Z�-�\��S���������W�rD�K������;W,�hz���+�LX:U�Uo1��P�̖�����{d��ƻ��2�	O7�lt�����Ox����/����BT,q�T��c޹/���4�§�l8���НU�!~bC�+�j��˙U�
��a p��/�l���,W�ָ�+� 	��PM���Xbu��&�'�gt�ɱ�VΖ���xl3����"�q-��	&��l���uΰ{�cS�Q��똿�Ӿ���F~��Qz��7���z�g� [���sg�rZ.e�.�Y���N{	 ��)륷��>s�Ro%�ڗ��]�^�n�z�X��b�b20�ʄ�E�����z�O=�A�!s�9����pfpi�@�Հ�� r�$7R����R
�]�܅�Q��Ʈ��%pa?w�8��[_�^`}����St�뜫� ����S�Z��=��9k������V�!%%�Fqj�-_�����p:}�SL߻@}�]�b��{�Zŝ��nڵ��q�B^']Lp�@�h˕,p�q�N�t�dތ��l �F�jԸ˲��1`<N��Q[.ӀOP�5��(*M�Dx���#�O�n�o�W�iO�U�K}��2h����F&�FFw�C-��u�������;�b���9�u�1`0��L��>�	�(�d�{y��h{hݳ����y~�zS�zU��sW�����HcG5& *��W���b\K$�J4ѨK"*�(��Lڤ����z��_U�y���y���߹߻��۩s��;��>��ϔ6�����d�}
���H���A��>�����X��`�Z���_D�}�fX�dr��#�0���+}���"�2H�hL�K���Y�u,��!F��ƕ����h@�_�}P'���|GrV�K�}/����:c��r�" ?OZ�Y�BP���R����o��%�o>�!���Am�� /}��.�ZX�ݺ;�a��G,����h�*>��(6�+;#/mCf���F�]��9X�!u�0�ԃf�*�W�];@��s8�B�-�����'���L��P<� ��my��`�[�Y���m%U��.�\ i>�я�?�]"��$劣㉇���'��/{�|�?}�����*�ts*u�G��&�,�`25��s�	�GZ^M'Ւ�P/�Yw�<n���*3x�3HK�GX rP��fGل���byy�C�� �>__��`���Y� �#dx�0�ut�����:�A����*Y!�{�=Y�ztB��]�=|�X���B�xɅ/��0ccՃp'K�z����k�{�A���6ôv�i�a�̕Z�T)�Ç���¾(�[^�)����ujXǛ�!
���������~�BwM�n�Z7%/�ҕ��a����,��Gx)I�J0֘�XF؇}�)�� �#�],q�`_J�D�ᒼ�|���W���8��4��Y||@�m��C+�E^�6Y���p����S �"�]�Jl�0�-\�E��>�7r��<[����;9B9]��CHc�apsQ�IsS�.�&�vz���b�;��D_�Ǿt�
�ȭ��b��TG�(jt�� ��.�ϰ����/�y�+b2msQ;����v�|���>����n�Y�c{e8ͪ�g��W�~�io�%"�+4��E�r��N�+��E��? �����ijހg�Cꬨ��TY)UM��?�2h�0�n:�q��4���y�9ܘh"6
�1���d�f؞:r��~�W��ѣe�]ւI�����#���Tkܫ}�I�AX�X�!��l��r]t��6�:�r�ny���e�r�0Q� �u��c�2}�f����W�z{RF�_���+3B� �HV��L"�sZ#;�|��~���kR��W_8�pǟ���뽇���,���BG�'�!���m�L8�˛Ij�ݷ;e�$��.پ�U���m��n�*èˢy��:���y�j�;��rOL,#�������B'E�Rڦqn��%�fa�w ���'�Z\��u�0�9yUW�n�2������]��q �j�`Ec��9]�X@�`�v����2��K׮č��<����U�e/׼ʅ��D�ʮ��]�����GG�����T���ػ���s��6oMn�@�7�P�z�*����k���W�3m�.��2:�$�g�}�����~qF	e�hl��X�P���Ġ��/�s�/"���D9}�s���˕�&�Z`Ak�Nw���^��˰4�,:���eǰ��َ������[{"�f���1�Ș��햺a3\�t�e/Mϸ�{#�!�{��u�|��ĸ]��2�;�}!�i!-���n@d����S/j�(i��w+�*+�~	�t�-�i�c8'���+����z���������c1���y"��qx�cg�+�Ǐr�p9y�ly���r���-.���$���π�Wi��R�5ʗ��א
�xuӮ<����s���4�2�]6�F���R��$�ӷa[�i�}�ߦ $�q`hHYt��*^<�]�f����}�K�Ɠ4����{�9ɾ�C�+tD�ܸL���!��Nr�䅛��o��r�:�� /��'��u�E=| �Q�w�{Ͷ]J�tT"h�n?u��?_֖lb����6_Z\��`����B�����l�fN��(�Q{�!W��mv��j�6^kP-�Ɛ��.����;	ri�g~�g���
��\ElJ桪��{��-�'�)w�yʚ�j˳/�o� �i�C�<Z.s����\b_ƥk�� 4&����sM����:��n�{��D�94�����:>H3���Ç�}hk��壑ր��,��$T�����0�ց(�v%S/�J�������3L����۵n��H�Ν+k�9�|��r����CW��Y��2} ����*�!U��z"�f�9�k��j�gx��z��ba�n}��s��񡺵:��g_�=>�Pg8��̛iv�-x�����`٣���ej+4XƬ�i�q��g�D���K��+E_��̓��0�[�E� ��������̙{}8��a�����s����9��.g����Ʒ<2����(\at�gEs���@4�i)��?^�����;0`yُ�7��Ȯ�� �pc"�������8Q����U/�߀�wQ&���o��j��W��u�g1Ǐ-��=��mwvЁ��n�C?x�L�f�9&������_�^˪�����<���P7/�6����	�k�l����@K����K�C�/�7�YgU�1=�V}y����Vw�[���˰�я��S=��Ą�`T�E�N�V[Ѭ�z�Z{N=û_�m�����ۋ|�k��B�?��r(�JL�\)�}��p^��Ξ.�O�D��U�9ͫ^G�3y�$�ο��$���}�;ʑ��+H!�3!��_��+R[v2�I"L;v����L�@�`cAyy�a�^$Gb��-_���P�m�~�J+����� ��	��Tש'�����	�M�4��8�4N�:�$�-R<�E:����.�a�>{��2�47��v�X(�i�$�jl#/�m�W��6PO>T"b"t�Ni6��ڲ�����P*rL�2�&��-o��<}�/�������I�_4 �M%b�_ڳw�@�0���O���{O�<�n.f��'>Q~�d�����@~���'���5�2�:��$���,v�~�V��=�t�^z�<��K����/����x5Ŀx�f��~	���[� �N�kN�;Q����~ J�]�*�b>d��5L����PnE|�L��7|���y����ܯr�������8��nB՝*��g8�t�C�i��o}����+���o�x�5.v�_3EĶs¸C%�J��6�u��"�8�m�&��m'��/���ŗJ�K%k��R����Oݟ���k�ݢ��:��r�P�rsO�*���гb	�6��@V4��Z�T�~ƕj[q�l�=={�1�q�����s?�s��ʅ%*�66��v%�?������w�Sw��,x�/�zyd�׾x�s�G�����E�B�vʽJc�܋ �
R)��@Y�I��`�(����CDs�A)�h�R$���S�J��{Y.7h)֌#X��0��@w����O�>U��ɔCls��-�U^��'�;KY��o��|����*C��W�&��%~a+<���r��G�9�����R��z"v��AuWe����~�_?m�V։NcX;>>>Ć���>��%�N����-���pC�/OdWi	e�U&��m+��U�;�5|��� �eC��C����L�S�?��?�����}eY</�ԏ?d��Ε׽�Ay��w���@F_I�JB��g���sϓ�v9{��������;�׽]��{����S�EQb�aѱ�@.���^6�TI��I#�^q�(��:wȼ�L�k����+�n��JK��bXW'}���h��\l������,&ѹ�!A)�OX���:t*�-W�y{��#�!u��Y?�j�4���0R������Ȇc�l䷧�?�����iy�E�ݕo�l<��c���u�eЁ�̓��y*&D!]�+��,T��Y{T����'��`0�At7DR��:n-EN�"�|������h���"��eq���r9ľ���J!z˃e������/3��s��+���2U�T�r����}��W���ʣo{{��O�w��@��R9���1؇c��:݄/�ϲ�zJy���j�7+� 䅀2�X�����<E��k�O ��K$�ѩV�J!P[��r��st��3tVz�Q����tF&� ����w�� ���O>^~�;�o�+�"\��)W���8�?�d	K ��[}9[��R�9� �=��Qu��\$峝�#�A:;"����n;�p�'+ٴ!�hñ����j*�[�Ҡpg��X������ڢDuO�/�����o=��J�2�Y[Z�9񥨹(
,)Pl�F��h���滩௨�* ����Q�����n~u�M��G�/��/���/�}�S���P*�"�3�z,� ����xac����o��R��GˋO}�얃"�#�tVHf�?^o��o��x��c����O~����rm���9�0˰��{._��mNf��/p�:,0��#�N� ���}��G�ܼ����"Ew�ɖx�G�}���(���,^[���'H��R����\9���{����K/���e���f�{;�+�_��vKݸ�\{m��b�{��]}0n��K�hC;�vf�-\4S�D�r�vg`�yWܽk u��%���B6>;�~dİ�Qq�Z�D,t�ӳR��t7^�B)2�/Q�	A25�.�p�=����c*<P���"{*����}��������r���${T��:Q^ϵiKW�_|�\�t��G�Rϗ�\������w�w���l��'>R�O��2l�
TR6�rm_Cj�	�$�f"�`cr��I�`sJ��O��0 @�N��t�CƼa�MU�~��s�Pec���7�8�����<Ĩ��������T.(�c Q^"D�An�����M�m <S"�~�T��l�����ƻ��M3��5l�,�z�%G9���u���SǏ��ulǛ})eٌ'���M�m܇�|
�
d�J����nW	L���~�Q'b"N��m8������>[�����_�诔ӧN����sL�\ق�MA=�{�[�¡ٹ����!x�w�G��Λ���Ēa�:y�{I�p 驏?���>�Py�����(o�?�����3_���PP��T`���i؇MV&���
�<nݘ�S��T��&�<:6³�y/������"��\g�tw���HM�����P� �U�"I��]�  vÒ�M&Z�+���7��s��t��鮞�0���6�s�cƉ�`|l{͎V�s*��r4ٹ�{뵻N��I79V��T�$��9���;
�"���B}�5n���5NB�w�R�!]�D����r�r�k���Ǹ�b���(�Oo��G\�F�D����!��}���������,�²<r��p�T���/�0�-(���j9�}	��9&u�H������3��7<ZN������ϱ�jy�=+W9�ӑAhw.��ߌS�O|���o?�ˁk�ؓƔ!$#��a�U}��xI�����L�(3\J��u_���T�������r�����Q��2�F�щ�� J:���HD(����~4K��ٶ]�nڍc=vS��}�9��:���
G��閺��Έ�%�_���.��2�d�X�~�IFD�~E�3Q+ڧ���fX�0�����=�*�13�#1pUO����z���P�����py��'�����~w�+���,z�y˛8�vo���*�s_*'9ox���T��^{����8�����ww^,�Pko�;5�t�*'�,XO������JN�7X��D��{O��������0�T�-+�$�}y�I �`*�d.:��p�m���e	�"�����˧^:_�g�<�,��ѵu ������|�+��D{����6���7��z�>m�������eZ��eD���s1Gd�c�$}� Tfo�o�LV�P��5
cO�*.%�PVJ�Dm�v�ڣ+e�2nW"�3l~I�[~T�(�tDr�wu�ӽ���Nr��;�>����������Ky���P^a��̜bE_O@��j�Uq��c����ڲt�Ry��,י�=t��6[cϟ/���\y�����پ�P/=���R��4���S\y|����tEE�PLe����HƦa-�^8_ƨ��������#G���'^g�u�P��Ti�����,{ş��/�=�)�!۔�%N�ó���
;;��x`J��H�D)���^�j���2TƲ��m�l�L?۸�f�4g��eq<6(K&q8|� ���Z�/�]�`ȑQ�cD�cI�m��ր�6�֣Q$� H����&�:��u���K��d�!ܤ�]�'�\AK�o����_�I����� Y'@��b-i�����sr�0HW�\)/.�䩻�r���������S/���@��*w�3��W��*���xq��O=E�&Fǡ�R�m7bQ�gΔ/\潝��[�	��@�ˤc�fZ��vO�-��MF�g��������֗`n���QaE�C�GϤ��e�tY�4���(��@�m��6��-!3�n��6�Ե�M���R�IħƗ�O��xE,�\y�[��=����7]�j�dV�,��d)�L� Yqu�Cy����WU��I�w۹Z���_�i�*%0uo��-����7�jG��.��|��ϕ��?Y����P.��ܸj��+� ҆�(�E�A    IDAT���gN��P� F@����l��<_��c2:V��\9��ܸ����7�7YhD7YŜ����s�8��H��YB|2��� ��-f�7�\//r"� ��g9]j_a�:�H�J�ݶ�9P|�R�*,���9l�:�УW`a\Nw/]tw����<��LFzx�B9�v�ֶ�0�}����[���]G�8^��.��h�2o��{2�6m�p'�ԺڝTJ����ws�[Zb��fp�����_2��E�xG� YH�Be%(��-��3n�FI�2
�Y�qK�3�a3�,��v��cY��o��<�������/�{ j|D�Zd&33�/�\�>�p�v���G_W^�_^���ǹB�Jyy��ԋ/�3�ȣ0�;�\ִ�"-"������(��DP��I�D�� �_�I���/�/Ҙȴ�Y$N.��s'�[sey�4�i�ʣ+��H�ZفAp��8�wA����͆w�U�-�.u�(%<��g��C�ݯW�_�E�T5���*;�J"���aX��{�`�����g�M7��g������s�v<+�.%Me8�K��=��3��qy�hYrÒ^1��5��PG������|}�xj���π�����o�x(�]3R�&��k�ȑ/Bi�.���+�)�꯳��g�=4���|\(���BL(.�RzՆ�A�oe��!��^���N�����?˼Ef�'���jlB���N���1*娓/+�Q�jV !P�P� �Qv7-��E�t4�.r�J�vt�p�wR�ak�^!��0��p�k�'=�}#�`#��ٙ�m�����b?����8�ߎʪ �
L����H@=�e�-c�7��K����9��� �=ٖ(?Q�5�ye�����?�+�V��?������/������K������\6���Y��s+�<o}�����,�\�x��]��B؄��2\:����{����8�
]f�HVa�S>_�-�)?����,���m�.���֛[������t����%j؜����*I����aGb ��n�!aM���dK�xm���p�2��8Vw�T^=)y�9�T	�ԥⰛ���������(9X�JOr!�s�4���-�,��_��Jܪ��CU��~�'p�g�8]T�Ja5�+m8K�JQR�ǧzt�g�Q1�8���>�ܽ�o�D��f���L9�BϷ������.���P��Y�d���{v��F8�
l��8M=R&���M��a3L ��%"�w�xY��-�ܩ���9�������{�l�E�~��O�i�]��4�#�cJ���Ò~���A�@��ZVb
BB;�xȦԡ���*{m�9�5Sݴ�@n��e�������}��3����zv�dKL��wQ��w+ ,�)w�}���J���BJ�3�(��
Z�A�[�K��V�\���"@b�F)��m����O�B�\
���}cg
����=Q����o�[�ϭ��Y�[ҼMj�x^�C/��j&��\8R��)�t��N�
�TX��8���D'����8ļJ�����7�ȦsP���ǿDIή8�D<���r)?�c�Z�ۑ��wU���Oص�4�x�*�OexS�El�j�ݎ������ٸl��㹣úmno�o��*�\�)�h7t�=v��䬻�J%5�ns�ͤ������4X6x��E&I��V��oL#fU������4��*n��X^gy|�\A�6��T����_�_����?�}(gO�.�؉�؛��6�U�a�;#u\F�� "a�e��]e�F�:�ԛK-���}�r�ˀ���
K��������� ��\�:�&d�
7g��bn���;�����U��;z��E|���N�
��'�/��4S�|�Jt���闝#�m�h���N���a��/����RӖ1萦:���o�D�8��u������E���YT$Wea�2�V�K����5n���]��7��)U��6J�ku��y�SDl�1{����h���r������nб�UlJ���'ʽG�!?g��[�=�L�;o�\$qQ'������y����4���*�S��Ơ_��_-�!���>����j�0{N�fC�A*�{��U��u4�d���?����RA�A�dī����a��#ᚁ�S��_�/q�vl��]w�2������#\�C�����>�����;�(�cc��½��hA4dO����UI@O
�G�@�:dIa�~-(�w%M%�<�T���wѲ�����&�3d�6�����J��O��[����N�����_����Q��F���q��{g&Ƽo|���?����E�;�I����=�����+>>5����F�o#�dס��^���� ����nܧ�;�_B�?��ߊ��D�t6����X*k��$�҅k E��7��j%�r	��u0/̱�K��Wa^�"&u4���?D$�"�m�"y�v0�TPwyQW�iƓHU���ŭ��zf:*�o#�v�$ ��O�DV�qC` ��!��>�8�5b����6I�һDp+ 5��OVl�������a�צ��n~�L�%E�R�'��&u�Ke>;T�3�Fn㛮�<s��/������gΜ������c������Q�ao���zZH���RVH��Fc������O��'�=���(��zjh�b�5�}'4��v=�~P���K��Mi{T8d���]R5|g	���j��������5t�����@�*���c��+����ddן}#�� )���$��m��k�y������T�'�X��[ [�[�e���i���	�L߼�O�����	��O�LO]������5l׸�3��|��T���g��X�W������?����q�i9z�K{R����'��?�٧�ɞ����ܕ�G�h2^ ���Q�`�Jn��d���kOU���d���!osIus�.�6�܇���/�t3�=u�f�q�!Ѵ�Sֺ8�S��e�LYj��!�^�����&�*���^J�' 2ܠ=��&r& 2^��l����[�5~G��V6���t�e���]}�9�F����'91�UV_�����^�&⎡Z9�2+�.���쮄�e�أ�NӼ���_�AӆKs�*���K�);C�XTw�f|]`+?ߔ1è'�mz��[?�ڷj���������������A�^��_䖣�h�6hn-;��g۹^��1��Oee�Z��O]�6f�S��?���xr�m�pZ5L��R��;K5��f���i��Y}�ػB�*9����e:���	}�$F2�h�և#�L�~
�q���!�1�(��[���J�Q:�UB%��D9d�z��aj}*<�/��u�6��2톷�}�DRY��S�j}2�fU�X�/�M�q�(s��Tc�_�r�az��ɿ?��]~���]���s�9�M�mj�gC�'�M	����v�\+Ry�lӫ����/"E`���ǯ�q�b��[g�~:�Ѽ|2�2Mu&��y�u�W<�s�����mʸ
Q�i	��#�a�t��4ܮp����\��D?�������0���WOs����nβ�u��8qmC�_��nW=a��{��͍�9�jaÞa��	7�(`K����j���E�/r�k�q3��Eh�68L9���값�e�z5!0�7Ӟ�U����O��=�Jaz@H�Å�:��L+�<E��V@s*��{�{=�m^��Zw�&�K������IŅ��]%q|�����=(�E�-R� jm���f>UYa�/w�+˨�#L����s�ѱ5Ww;��ѠYN6�2~��]�4�Ѫ��`ڪ��^�L3�kX�Ϩ(f���x�bBX��|v�Z����ԭ��Y�xQoF\� �ET����Ut�rd%�?+#|����&� W�A�_�N��K7����4��^�2LX���Rtچ���a��u.�T��3~WB�c�l�k��9.I��ӓ醷�,�z�!�,z��a#r��{���i6���0�M�[�6�L�����X���c���6��v��H����8ER_݅�0�5A���i�}�P��-����Tְ�"ւd�H1�ʤ	�@�_3?=ʙq����`�K	s�gx�צ��*өY�*�%�����	kqj��%�8d㛶w�YW��uO����7i��g\���n4�x����7�y�����E��dˊĎ�Z�
�d1��e���F�rZ�N��V){M��n�~������~��!I����	��cG$�m#���,O�j��Զ��^?۳��>t�׺ny��j�������<P��\,�3X�l]Av�o������w�K����x=�U�~Z���O�aURݍ�]��W@��5�z?	hv�[;� 2���0;��������h˓ygw��l�:f���i���?��iԑS�֞�|��nYu����ؼ����9��.�;B�=��{��#w��l��A����W΢ns̤O���l��Ӏϴ� �*@������5L�͘]ڤWӼݿ��2�l���DTA�n�'�i��=���O�~�K&�R_+��ܽ�<*�J���O##_ޡF�%V�L����9a�{F;�����t�������p
��̷�g�M=�(s���i�k�$[�9�-�s���޿�G�zJ��n ��Yz_@G�q}c=��d���D6��}�>���ަ���N{�F�z��0�Gu�#O"~���Ks=����Mo0��t�fo�ʹ��z*�U�ƣQӬ��􅁝�v�~���2��oX|{m�{�G�D��2�o<�-^]D�?�q�2�w�aP�7r3pX�!2��^�
V9фb�%xxL�'��*����t��v6��&P��<X�eG����Ul�x�=��|��(�e�X��W�u���������&Ŏ0w�A�Y��0���D����L���MЮ���X�z�q��Td�)��C�H��E?tpHa�k���Q���
��$��4#��tLCjN�F��p���k�;Ŷ��#��ͱ�q��|H b�k2��_��V��-��6`g�t3\�u����,�q�Ӛ�f����f���^�$�ݦ�n;C�mm��,}�j3�f�����6m�m7;�_�׬'�:_=?�I�����^"r�g�A�iH�UN,�_]j.r��s���Sn6v��ٌ���w�I��j\wY	�Qx��-�tEI�_��T�O� p/섉����l$ː�zi��|L�0.�QO�;�2���
�n�1�{�cJ͇�u�IWU�q�� ;T�	wEf9vh,��Qw����6�y3^��()�n�XuO<ݸX8*��Ȳ���!D��-¸hf�m7�)��q�46�+���*�3�����rM�]T?ջ��(�p�9����@�֩qO�׊1EV$ۚ���n�3���~ o B�8����L��Ӟ��l�	t�U5(Z�����ʙ�fy��2�H���8�ӎ�Z��܆׼��`X�Y6�e�S$g:i�-�-4믞f���a�n��mޙ�e�J���
'D�j������M��9��[�3��K7�	(v ���r�?�S(�h`�a C�.�36��į�SUy5�J#�>u��4c�e�"��VM3�l8��'����Fna����g޵�k:�Qӣ$4��1n6�øď�&���$�
�KMK���*��y�Y.�fU_��Q4Dh�l�q�WF�яol�;]:������xN��6B����V�.�zv��I�)	2Y~��l�?���1Ľ$�1b	�V�|c»1	3���L'���>�e���;��} ��Z�X���\.ͯ<K���Ͼ���,Ö+o���ڇ7�7��F�i��=�5���V�M`�/��W@�n��+�J�0*�UO?�M�C�C��/_�?)�e�Mez7�g�,�nqu���ߦ�_�������uw
�����Ջ=馞��D���,QVt���u0��:��I�gx�2L/==Q�^�U�d���k�s���w��W�^���:@��>��������,�x>�������W��=v-�Ҝ�H$Ю��T��n�})Ag�A�#T�g7 �f��;��Yw�A$FS��=�n�W����4#�.�^"{�4�����K�g��Tփ/�a@�{�O�f���Q��mq'��5t�0ӱQٞ	�-����i�/˄~��U1�tW�I�-���ԍ���gߔ����b��Ec<��}sbj�����0�N-���q(*KwTZ t��W�h�[���Ġ����z��O�q�_?�2�l�A�tϴ�[s��b�����kˮ�/���ɊDZ����]y]hD��mm|Y�ɰ��W�.����5��a�M��+�U���8��Y�{?7�΅�?�Fn6r��l��s��f��=lx��wSY/do� ���e�l� L��f�oU�{��V����8Mok�k�8:'Rg�6O�e~鿗^�!��j��d�uJ
�S{4tJ?
����� Z��1�ƿ��G���\ȴ���0�eu�U��G[~��5�>�[{��8��Un���,����"ޕr�_3�W����'O�����������to�Ѡ�B��=+�]�� �� ��4jO��[�q2��3?�f���洧�q��;����1���#�e���龛��o�i�w��nY�����-w�@���rKLZXePØ��*a�s��3~�.˓q�˯�O'㙗��i����f�ϝ;�̾w�����	��kE��k��
|�!� w0m���+IY��-x*+$���<Zq�3^\���t3ͭj�����3��gg��������j�u��#Ы��8����֫Ъ������QM6Ds�	s���u"� �T�N��{�Y��Ȭ{�k��W�����0�����ޱ.�^��4�|jiq�WW���^����=����>=�������{��Y��da�SY��J�_�מH�9��f�V�٪������3�v��~����2L��|�<&��S�i������-|�g�A=����5*��*�}�$�L�6���Dp�2n�SOx���L;�d:�J�ZV�<���'s��WVxY�(���6�yw�x �n�0�����;l�w��D�2nV����;�H�;������Z��&+Q��i'@Ե[�l����8��k�e��lt�i6|�O�uw�A��6�f�QO�O��=�S*�Ր����+O�k�]�Z���&�֎�g{�j��$�l9U�%^��캙��l\�х�W7\�Q_�H{���	s�Y�����[�M?e��؋�'M�����&��ݕ-�7rS#A6����}��\qW;(�����l�[D��$��,�.z�1,_V8�i�_�|�_���5�[�zz����"z�g�5t?����k�w�oöf�ߦߖ!��:�~��b��2d<�7�[�M{�e8�������l�}�B�ޓN�G)�hutz�����n��ۺ�
�`[=t�3o?��s�7�ή��sQ���~Y!����$�}��[ȶ���Z.g߬�ƞ�[��Q�[,w���}�[��j�v�JiDlU�=�E�گ�T����|}����i��km���-��]�i�!U�n�|!5��ȓ<�$x��"6{7�v��*���?w�S�Q�-B{@AQ�����f�x\b���)�t�7�Flg뎱aʓ���Eks��{K��BZI�Ys[�Y��E��2N��፟ȩ�ٯ��m~�� �a3�ަ�_k�<�]=�����=��� �_�u�uk�3n�հ"o *��H���4U�f�¡��u�Z?���7h�=<����|�e�2��m?�p���f��m���2�]�}#w��:�.��Ӏg.��*���r����0{���/+�{=S\�kz-u��ߡ�ׄ�� �5�ifGJ��?�ճ�GW�S"�OC�~Y]��sF��Ou�;jOe�_��q-C���h^R��"Y�$!�w�jm�ȓcWEǀ���`��0E�!BZTR�FV�<�=ͻ�����~�nʷU�J�ئ#�����Qݻʹ��ܼ����ZX^"Sa0�M�����ّ��M���۝T�I}0��(b6�'Rd��W*Py�;���|�o�t��Ӟ髧�z�k��kn�kӕ@��#ߎ�h�3����=t�&
G���Mwqƻ�Q[����q�K\I?uݼP%��Yx�:̼ⱉ��5�q��-����w�����=�ek�{}��5�E�+�K�LQBB'��T�b��    IDAT��W��)J�t��a��=���6?X	�^>]<ä��&��_��i�#��8�9/�7L�aڸ�1g�g��UڝhQ�0;x��7���a�b��q���e�v��j~�
)�69�ۺf9uKs�5J�u�C���ԭ��7�*5�=�@r_���<Y����� 2��O~�|�����!d�M.����u�;���� AQ;z`e����ʳL.��ig>�i�u�<3�z���n�{�=U��v�6��}?��13�uK�L��$�fy�rf�W����</�n�ӭ+,�=�=�gҬ����n�+��B�@m�V�i�I�7[�\;Zys-�t�FW�3�L�يe��̳"��=mȦ�w�� ��d�=��2�LW�H�yj�<#\�-�,���E�T7b��bχt��#巜���s��o8cd����Ġ�,��R��*#:�mq߉&K�Of�6��^8�~�Qe��}h��ݩ �#_k{�L!��ʔ�)e��ŝ�H�E�M;^G���ޱn�*�h��Ӱ�	��?w����V�G��g�c<���EI\b4:��L�K8R��g��ݥnsParb�[1��Z�������A$��U{ �^��'�5�t�-���8*��LO��m�̣�����3�;�J����S�3H�߽}�3M�����Z�#,���_s�1ӌ<��+P�z�I�H���!<1X��b�~v��|��-ի���9�n��;������1J�����Nv϶�fE+8'�@EW��uo�����=U�����=-wԓ���Y����y�n6��=���[�ߍL4�v�z�g����n�NSߌ�.��&G:�~��~�m:m��%�h���sϸ������[�iʘ����I8݈w�m*����L/�;�u��}gg.&�y�6���[��u��-c�ݔ�6�)d�Փ�nF]e�l�Aզi�L#�����<N{���n��,�ni[�TmY�m�8�e��O=㥮{~�z��7˒a���ކ�p����n���f�Գùx�{�B<�kO�K+�vK�u�7�f�,���
-�@^Y�M��`Da�{3�Gg��ߠ�J��e:��ֆ��9Û^旺n��n�{k6ܗ������gڷw���zp��x�յ@��n���.p6zv+�vsҚDG�b\�F�^ڤ��qSE=;Xf����'��Ӎ���CA��e�fK��KoY������U�������p{�w8��E܆���`��˟�r�z�M�
��n�m�*���	����i����2�Aw�;���պe�>�_L^6�z��i�g��~�M�dz�iΰ�[��F�z.��z��{�sl��(
\�ۋ/"�^�b�G=��G���l�ѣ �C<:*��3|l�,��\�"�*$��z�`�X���7��x�q���5L�֚�8m�m�/�l'6��2=���񮤢�u�ޖ+�Gܻ�؆������-�H�{�5�6ˮ�O�yd��=�Ͱ�u3|ύb�(�̸���'N�oO"\���I\q������:�k8��/���,������
���a'$^Gfa��<Se�'`�-èO�a4���n�t�4RL?�gx�v�F�KUm��&-�[�^�;�i�i��:�W�5�o/m<��0J�D����<������"ͮ���[�#���q�r4�a�<nܨ+��}�˼�y��>=��=<���-�l��. �������1��mʱ��@j�WP���w�~-r�/+��L�Y�4'�ɰ��f�m�~m���p��J{�մ�qSe>��Ꙗ�6�iti��ƕ27YGr�g���tul�O��[����]{}��Բꖓ��]���~v�]?���&i��7y�t��m��w.aڙ���'�3�n�;�����
��#�w�l���g�l	p��J]��zAO��f�� Q��ůV�/U�-�f�VY�T�P�3|����7�N�_�q5g|��9�͸�e�2��K�0�t7M��k�2\�����`m�����o�hnå�n'��kuˬ�1^��a#�9����X>�M��/n���=.6�"�8z(Q"'�۩,��9sWܽk��2׍L��e�d�FdFq��fȹ-[�z���]�X�p�,��Qw�*�����ӿ#i�m���2�id�hT�����|0f�W�Q�Y�^i�ѽ'�Q��t�e�p�QJ?�CM%�u��xY�t�Mw[���W:�|5e��{���OЌ�z��G��=ӳ�!m�k������"t}[�����k�q�[fW�C�܎E>�ޟ��*��Nպ�Ӭ_��ά_����=��O�i�kW�g�p�~�=�w)�H��R��}��F�rd�3��gg���ʶ#���D�����L�g2�G��+4�����0k<���ӽ ���O���D9��rAG�ۓ8�F��~w��M�y�A����K��6��Q��݁�V`d%�0VZ5<��g�3G{-�&u�MՆ�M{���n~�iؓ�*�ɖ3�o���~F�>�^c�{��i��M�L����'z������4Y�V7���Q���42^��h�n�4z�3���Twۢ�����ק�y1-ٓ���a^;H�f����FnX� �vS�h��?�k�kX�Y ��~[)����m��j����id2�`z��N�_v�to�[��t�\9,��_��q�4�U���j�Y��ph�N�֭5g�t2�z�k"��;�x?�3G"^�P�|ϴ񏉦q�s�fN$��m�m쒾��o���2 �L��`S�*�ʡX�D���pP�D{��=�5n��j7��~�3�t�3�tO��z�%�ʔz��x�z/�@����3�i�{��@:�q�+�n��-�3ʹ�H�[�4�f���fôj0\����a��+-a��%�HBҦ=�;�����b�T����\RY7�D��������������uvj�r�����:{Q"wL$1Ǎ��f��J�f�iO�hn��9������z�@&ͦ�*�2^��a�r2�f��z���ץ�i[�Vq��gm�i�����2�F�c��/�Id8�/�Ro��*����ZQ�t�,G�A��a�H�t���(o'H�?�TE���p}M��Uԉ�׷���?�FnVע��1[��f_�D��l%��d�2��,��7��Jd�Z�K���6�u�������܌�j�~9F�� \�z�x���ȇ��꣓����i�X�t�Uδ���a�׏��{2?�T��nm�Z����F��bF<��Ong^'�+oRw����6�ʜ={o���	&FK����Y
V��ʒǧ&gx�Έ���1*a���2`vTwx�A}-���2?�TO��t�J��H��3���;Xh8��f@��Xh�$��<��Ꞅ�x�c����:g�U:[U��^���"m��(ʟ{҇�q�$i�ӮDV��7yP�Gj�sNhp��/ab�=&���IbO�o�n��gE���ߠ��>��-_z Be���򧍓���=�$d(5�H�ig&�˸�Ty9�f����9_QN��k �P��3(�\[Y.ss3e��R��ˋ��G�����́�X.^'��|˷�?�_���
B{�(8>�$�ն������/���g��BL����"��yx@�R�N�\MI��܊"�e�N�^�.�:RĦ�zv$�]런�#��.�U-�zp��R��_;��٪^x5�w����Ӊ0]�v���#�|)r5�l���8}�5\~g"�b����G+
eST�'�VWI�SUJC�p�@
���HD* )�x� ���� vT������c��'�b�d�
o�;J������Җ�$�v��\��y�^N�{��ݟ��r����Ʒ���Z�g���ۙ��賵�X�\}��M��H[�?C������~�7���;��<��3��C���%�����"8��6"Ј��DT@���P��H�b����L��4-B;B�
�Jd.��G���X��[=��ꔐ��#3�4(�%(��a�_J[A\̹�p=FDPj����H���r}/EXB]6��xfud��E�j��G�x�2UT��X�A��7��n6z�3N{�~f����޵1���W�W�B{�ڣN33�m�J98;Wn޸�9U�\^ �7���گ.����<��7��Rϡ½-Q�'?��e� �mh�^�+C������,��
^���[������ce�ȁ�|���?���W�cÕ�1oG�d�qU��傲p������:�fWg�1�޵%�G� }�g��lͫg¹�h�F7L�ӯ��!�~]v�e��#ZO5�^��S���w_�ϫ()9v�X���ꐭ����`�7r��e�Ҏ���C��#��7͂����S@:+�[y�k+�@ɰi���q�EH�D��=M^C-�ٱ7��9�������R�n)0/_�P&aU�a�W�ڟ/G�,���@�Q(�X����z�*� \-˜�C�A���g׸`���h��5̲7 �ƭ����{�3��w������r��8��d�yG�/�o�*e9G@~_;Du ����o��� {e�R�@�h&�����'�G�5���7m�O�F���_m�l�q�)�!��1���F��N��B�l��������\�w'}_����������$������G�`$�L�F�2���-��#���h�
0+�{ �:� �v�!|�����>׹���ި�5�y���s�9��Ux���J�k�W
Ѓ績k�|�w��������׃��v�
H3�q�	�h9r��L"���%�����8_&� 7�Q�����́p�E?u�^�|
~��B���J6�*����4�NԵ�@�pՁs,���z
gU�b���֝�f݅M��]2�����_d�D���i��e��-ä.��ٷ�5���_~�r��щC�N�6+���=:>�q=��9�l��y#ޥ��y��Y���n�VJ-"��2\�����}*�q�*�@�|)�ʗnu�[D�0ye��0It�͛ 0�~�W~e����r�� �+\�?_�^�ä�~yy�LN�����ū���	�ݙ�aX�_�l��
H�y�3X�i؏�7.�q���^)K7��[<lt��da?|����{cR\�+���X),�p����p�}�jV���]������Cs�^=үI�~��ԺB��Ʃ�4�Î�e4�NI8Uۖ�v �;q�D��U�2�i��H�2� �wQ���/���wY��q���o@�W��V-)��[� DB�.�Jo)PV�F��dD�g8�2l�Y"�@k�䷕��_K�"��[����_*����ჇA��r`�`y�����q�M.i��ˡ�sP��6�a�౫:�/߲�K$¼��Z��)K�܌nL0�X}���t��\�l��ó����ꤏ�����e�NW[�"P Q :YH�QN��ȦN�D��	�M�
�|;'U�*탰�=ag��+͉�3R�'�[�^(Kg0_��{��c�VWE�*�
mż|�Z�����ͯ�X�����7֜Q�ܾ�><�-�D �t\j��������k�ʉl�J����D����#eowUk��,���QB�%[Q��>6֟������[ʛ����	w!�'U�2�E���;EF%¾, ��ZE��X�>�V�ɩq�?T���4(�fsk	^���n0�^.�`T���T���(������J�VaM��� G�B���+eb��:���L��ӫ�k�^�� `����#�^�nP�32`�|y����R�P�	�w�{;n�)�1jG�B�)Ͱ��+ݮ�M�]dh�ɱ؆B۫-��rk���~�j���'w���}/�/�]ʷ�l���^�5�j"����* ���q�̊Z)�KU&��>��Ͱ��d�Z��5|� ����N�$�ȑ#�sD	9�,�d,��������<W����,��+י��bbe�7���2A�SIDuK�e>zll�k X����v/��$�-�X:̱=<�F<�G>;�oxd�,�|���C����W*7�/��).��^�%�����Ab�$�� �R�	���K�΅�=��������O�M�����m�,��(}�x	�l?��	�#/�vݢ�;��a"@'����o�Éz� 6�nӔ����	=���Lp}_�}������u�n3���8�r+G����iq��ʷe�0�%b'�w�%�N��_��]�"�i~)��q�A)ȱcG�&qR����K��`�u_����Ώ� �*��X*d�1���< ��fw�1�ff�=�,�CJ7_+�P���_����cz�S%���\ER�� K���,��vbb::���f��*z��Dy��3���.��(߶����Vοr��Xܠ� -�.���9ne�E��x �λBgr@I>��6G)�U�_��#�}5ؑJ�T?�;��4���ILG��໵�YK�	�1T��<R�9Gn���m�.��U>��v���ܣ�ܨ�bi�.-l�,��������e�,`���+ ��'�&�G�L =�t��;�2h����b���PaYCj�p��bʷ}۷����{���O���z�I�*7v�ƅ� �K�  �敠֛KP�eq�2io�C#1Y�	o�L\����,ȸ84�����3����k��.W�!����]"��x��2[<^>���r�)�p�K�{(�ty��O�����Ay�%��	D�W��,Ӂ&�8Kt4���I��� K�D6F�4����p�3L~&(r�%�U6ݴ�T�q���Q�j�I�쬟��B9s�yF�ҥ�V�B�6�%���T�zcD���~7�xR����;����5��m����Hs���ƌx�V��~����0�����wѝ����}wy����C�'�]���ϰ�a�.�27;Ų;T1����-X	d��S��˅K@d�h�B�^,�K���k��LM��	5�Z9vN�'�2Y����30cS���	�1�
�W
���������˗��O-�_\�,o|���#?�����?\~闞$}�X;������M�׿��
�p�e��]�1��ا�����=H��P����v�&��4�t����6��{/��jbb$ؓ�����c�������;��ω�R����5�غo᰿�E��Z�� �պ��
��h��WO������ęu�y�zH8(+���޾���|���E�9� �6����|q�I��R�m&��K��U�����}��O,�l<�LM�Drb	ȑqyB��$4
��Mf���,)S��U`���H9��e�ztd�:2�y�tf���rz{�{˵��'˥k����ϗ�O�����~�)��{ϗ��?_�|��r��[�|>d�#�[g ԃ�bP�@�mR���RdV	����?�t�v��to�N�ȡ'çn���/:�fG`�\�9~��Ёٙ�龗ڽK����"���6��GJ��F�xR-�8+�%
��v�|\_�d�������^�5�F~�b�.J�=��"�
��р��n!~��^`�������o��߈�׮]e�u%�k]A\a�bhg'��B��SS6�|y��ϗ����@��P�u���ˡ[�c�����/�O��2;��n���V��C��3� �#�����K�0l�ְ��B����ÓX��?�X.^�h�F^�j9��d���PN�:Px�x���|-���)��jm��I^o���<�TVJˊ�C.�+��K8���O�JJ�07��F�N��btP�^۴v��sd{ն��:e9��ٮ.�u�p۫�o}+,���q������=]jw��Ŗ�]��9�$�r��=%��\[c���*H� !nx�^�V�Ъ�c{fcO~2��4�:H6��-[��tӬLԕ�{�9�$�����������A�X��K��^�>Ϟ��@�nݼP.n�օ��z�A<�ݤ?��>�b���mxk�q.E�j*C�Bg��iD
���Q�Q��%�5�F�xG�D��sK!�^����F <bL'�k[A��M�-�_x��tu�����v�E��嫿�]�G~������b���v(��P16H$L�������4'��`<����@���v5|�W�$�팧ҽ3�8��O���1��/����O?�4���&DV-.$l�    IDAT7�Qw��Bn��!����6�׷��s{)��8����%� ����Nܤ]#s^I��w� +@ԿҲD��<��I6yE��[dB#*�0������|�W�BT�P��Ef�B^�$�}쭏��}�/S�C��rm�O�[\�R�ͯm\�dM`?��k�W���4���H����Z k��3T�m��^+�ť 9�_�ޡ�%S��L[�md��/ D�Ed���|��	��&c~����jϢ�y�b�
s�f�<�j��_|��9�@y��)/�|�|�w~My����G>�I�����h��r�nHV��I�Wa���"Q$�� �A��h�!��/ʁ���eG��l����0�v�hGe�T5C �-L�9U	L,L5!� ��Y�gy�u�,o`!i�w0�{����)�V)����{����x߀2�Z�Ae�+@�Lu3�a��HѦ��җ���"�R����d	��;����W�ǿ\���7�^���<�����Di��IDv�`]���\������TtrJ�(֣��O��D�I\�2�j)�TR�ӱ���p:�Fa��E� �,;WC�`ǕOg�`�Ō��4�PpxP|@=Ţ��`��W~�V=	>5�uc婧?K�b��C��B����=R~�_�kF�U:�WaGY�B��(����Ŭ�*�M��������n����Źb{�v�i�������ؐ�z�¤Y='���#���xrr����ȹ����l�r�=��мڕ~ƦG��:$g��Z�@�[��_tW�p��pȬ���6�65�(���I>�}�(��Y���������+ސ����(tc�=�P�!�|�������XLaG�6K��K���@Mi�\����mv����bI�JLR4�Qc�� �e��ENp�ӄi��CL0ch��[��~@�qS�����(�<����a�S<��j��	�㾧<��2��������b�|�����n��-,��Ú��P�#���[��&�3$n�iɭ94�խ�TY,���Tݶ�.Zk�^�t	q���[�u�vM�	Oɢ!��ms˦���go�/����B3~J���ۊ�ږr+��u �9U�ڳ����Tm���N 0� �z�F�ڊ���1{�,�C�>���'�xQH͖It��H9�#�^�Zo,/]`���<?0 �+�L#�'�v���7��3�dug���iT�,ӆ�8��Hi��r{�4�> 9�:t��A��!6������ �=Ӭr��3�З����3��3���}��{���CgCl69����+�����}nn��c2d�9��v@$O
CD.1��N�8�Dp�+��K���l�A����3�4�ܵ�\���M�Cح��.j_�m�ԁ&�˭�e�-����.��Bν�[������+�� ��B�X5h�תL'(�'�M�ೕ�L��</��	�x���]����!b�q�z�7aC�K+,��h�[�_)����ي���r-�C(#�U��.���1��T4� �e	��[Az(R�.����\�R]`E�.��4H��q�E7y�j�+��A��l�f;�Y�|�ۊ��cL�op>�$�>T�y�Y��\�?���ןe$�����|�ϰ�q����Cl����Z+���V-azM5ipy�:_�A�{R�����5>�̿l�a�)�S��N�$_dv$"��!N�C�&�Vc�s����c��L�븳���履�[��kkt*�?P�A��Y��l�Y�;�m���G
�)�×�u��={_9{�Y��c���D}���[�!�[������^ ٖ
s�r�� �Jt��a^�`�]�`�%V���n�YCN�T
�������]��9(�Q�8yb�r��lh� ����q���g]�f�<�@��Nv�z�_D�93�\v�i�V�)�jy�u���˧>����������{��]��O�83ð)�#�&:L�6	�
�7H�c1P��S�Vm��aj�D�Ԡ=�S��6V��e9c��+��`rw}_�mRtFI�⿡���IVo�T�� k����*K���	���H��2�n��6%����
�c� ��~�`�{������C_em���|���ɣ����x����]-Ǐ��� �A^�^Y�H�r<�emyj�r_�����&���A�`��g��J#�&��Ll�E�>?|�<�0����l�9��d&a��H+�;��/U��}Q�1)�n����r�=����R�EʽȹN�K�^~�W~�E��r�����g�/�FD�u��1��G
U�O	��	e�~�)�A�У�$���� ~v��U5��K�V;9 [��&�@I`�V�bK6f��N2A�z0��j�����2T�;�(Ȗ��ٹ�J��Wi�a/e�2n@7�v�A�o^{7�n���m��w��]��q���ny��s�M��͛��~]d���ؔ�ؓ�����Ԙ}%"�Ag����xk��D�Q/��	����@��5 - "�<�,!�'�0;O�2�2���Wʺ���A�Aٙ��\��b��F�D�׺���;�?�����'O���y�N�	������g��\���O�/{�1ح�����l������BS�6"J�P�%��0���ٹ�[\/���h�ʥ_�U��/�Q����OGm�%y?�q=���V`wvNLL���
��j?�=�6��6>��uxt�R�b�ZY�1�L�����iΊJ�����_]d ���gxӏs�l��a���a�+��?��7�7�K�.���W��D3l�f+L��6�巼|��K[�� 0+�na-HP�An��A
��v˪�j��ǐT�pCl��)����J�n˜f�7G�9D}-����H��������zZv�1S�*�X�5c.�PQ�/<:ʊ&,#�>�F�*��:
W)'˛�t�|^�{U�?��)���}����);{�)���F��8Ƥ��������d8yn�t�m���*[8&ǘlW)m���VEےL?�>q�6O3�ڎ��z#����ro�d�2!H�7�˽>19�@��[2BK�l �Df+����T@�tϲ�=�t��i� 5�圣���ه�._�o��U'�L8���q�E�tj�ʱ�ocY�ɛ[W9�H'�7P��e��|TJ-eID�M('����[ 7�?1q�L�jx��Q����9���|�uB�Ȧ���4��h'"q�l���G�iE���0�\2��Od�����l���&�+�`���3�:u� ��O���K�g˻������?^>��%��
�?�.���#�u"������L۔Q�"H��"L��8�X�g�<�;d'�h��,!���숬�5��?]�1+���Ʃ�W�F�U�U�c�[_[�➍z�����È���,�3s C��9j���z��k/'�256?��ᡃ�����?��������Œ�R MI���H��1�ZE|6��P�FL��s����2�]O�ț���~%�0%��h :.,�v�!�&�P�9���a�Ρ����|�o\"�u�27�-r��$�I��ᝡہ\�h�\	�"� 4�p�rJ夤"�R!E��`;:���Y����p�C�3�����#�R������Hy��G����-��g˯���('��|� �#�#�l�+�9w�lO���C��\�T���Iwu�@"������ҏ��Re���4�𖧆�hB��Ǧ�/��?���e��*e�d�}��%Ûc�l]\ZdQgh��tH-X4J�:[ɬx">5��GEDvT�	�~�|4�p�p� �,�z�;��w�}����G�S,\�����?8;�􁳍����!6(�k�8R�^������HVDn��lَ*�ˋo������,[��{7�/�l~��+PQO�ߢqq�L�4��9 �@9��v)�&���v�<e	lt	��nd�"�Hb'=��D�ƗU[^�IǞ���eo���R9{��r���m_>\>����t\&ǫ�����_G:$$�rұ,�Lě��S"o����v�uwس9EX)w}"����ϭ���2�(��Gۻiz\�y��7��^f�X\��� o ʑLɟT�r�����Rɯ�H*U�X��J$�J%)W�"�P�%�e�%SV��bDi;I(�@"@ �%,vg/��s��f�<���}=�~3+���y�~߾��ӧO�>�M��^/�v�l�;����N�ug�;.�C�=�<rnfn
V���2�`>,+oq|���o�S��is Lt ����fD��}za!V�V�n6O�	��Y����[�h#�&�y�[�]��<�6C�G) P��w�GG<�*2�=��x���恊Р�O�@�r"�}LdQQu���@(�@�J����[h 2A�Go��6(T$�8Ÿ��9׮�-��!��<��F֜��*r���Pa��%��ҽ2tO�t�?`	R���5(<�O�m��������	;�|��OQ�s��=Ӽ���L!�调�0l�_;�4�N�{9eU6�N�&�r��A�Ei�il۳t����=	�,�����ᅭ��y�fL*��g�[7�&�ve(�>r7�m����oݞ��_�=y��=o@�1H9kﻣ"�X{ؓZ���Q��}2�^��ȓ��F�?��⥋ͯ����7�-���D�}%�����NN�Dd�-a��6,ɶ,|�{Qw=�z(�,�|-lX���EU($ϼ���-��[��a�#���\4�����8���
����.�Pw��N�ha��Q��6�ґ}:��OE��҈�R��J�Ο?����u&��P�]nn߼QXf�r�?����^C��B��<�#TN$�X��uځl�X��Du�~�v~k#�滶�8n�H�L'ڟ�E�dh�IVlmK;��R�c3�<G�c!�����ѱ���	xl7q�"(�h�v
$���D�9���`�2L0� N�6�x6�1����ͩ3�l���|�cO7�}�2�bV�6���{�E}�j��M(8�W��(��E�Z^{���Ԏ��!���@�eA��	�ڃ@�!\�)�r9�t�?'�P�-v��A��;�Zw�GAN�[	�7uDh*��@��HKG�C�$�K�и���<���vXҢ�v�P�%ٛ1�?yd�fd١,7o�`)�BP�˗?м��nsE�S�G�� ]�����Oތ �UF���Wʺb���SW�;���*oψU�r��,:(u��P�@X����~�X���";la(��#ͱ�����橱����m<������v-"V�X�w�8)p �J� �t	�� �~��,t�8����왳h�-�󆼝�a�r�Qf�U�����/��x��2������Y\hΜ>	�w�!_k�o.d�SdJ��)�cL��/�%#��l��~���8�A)��.��qO�����K�]�Q��r�4)
�v4��è�dމ�������K�c�騒���,�ad��],�.4o��Լ��+4��|ꙟ@\�d����`�9�C�k�N��v�T�إp��X?M�����^��s{�eJ��[8��H\�3���<Ta��{RW����0�Bp�]Wwzjj�=��r{�ܹS�� r�bpϸ.�R8�,���r�n��}מ��]�H��t[ʪ�H-��N[����� �V!�qa+XB���H��,γ�`��.��;�B	I^]Ʉ�>�urj�F8�t6�~��`�%��f����; �c��P�R'T\���F79�O��&�j ���K��t��u�CV����+O����� �n�����:���������&@��S�2k��.�9����=�D��}��?��\�4È�X��g�h���w`=v��'O7�,,�09��pb@�\��{ �m�[>M�A!FR|�=Qd(�3�H�J����㢻�p�3&���i(�v�8u�D�ХL�K���s+.X�#��� � s,�F]��eK0F8Df����3g�R��8[�اPD7VD���"V,�
�����6�t�h���z ���~�s���.E e�#�@�[��i"� *�Y �P%�(ťLPKQF���(ϩtF^��E���s�߆�B��6*S��vq�C)Ï��l�*utW��9�;�T� :�?� ���v"(7��23
8y �B4��x�?i���n��eP"۲ƙ*� ?����ls�6#�D��gcʹU
1���5�T����=��o�y�Hem���2;'��3�5Ri;��̢���s���T��⋝Ev��#��t�g��Q5:Jav�)>α��H2�,#��q!5�EX+��n.jԀ���E�|7��J��|+�8щa�s��_�p���[��� ����w�fc�V�`I�*�i����9���4>��{�ܹ�w��|b|�Oā�kk���e�1#���AY)����Dh��"�R�Clޣ��bv��<�vG�<�n�ߋ�Zg���OJ	B0B!���F�d��S$'t
�-�-/��Ɏx�2�_��:2�A��ANB-���6�Bn�����D\��2�n����.�?��E�9@l�[7��G��$x��ӟ�bt����DsJ�����@@�h�� âǖM�D�a�>(C�=R�3bL�����6 �N� ��&=M�~7��{��C�C�2^�� ���ab��U��,�#�6�?3�s׍TT���A�">*�p	�G������˾� *,M1�3��B�-�JKm�jzuR�P)4y���a�SyT����OY��Ő&~�0mt�B-V+	�>��&:s�@�6v�F[��03�����2Ɗ�"G1{.�;�pz���a����˨K;ʘ�dގn����h�Kw�i���u1}�vd�7p�#v@�}�+I�m�ӧXu�И�ixD6��:�.t�+]��Q<"���6(n�"������X +��P��6��ɰ��nCGÙfĜA}�s��|��*��y;,r�*ɀ=��4�i��md��6�G��eؖ�s�
�����	��ὧ�NCV�:�/*$M�3]<�`X�`�����*�pQ,[��ٜ�Dը�ҋ����T�z�伌1Z���Pa�O�Ex~�:A˦�iB��N�B���O]H����	��zz�6_�o8�������Ia���Ňn�����z�6eW��ZPT�m�)
ʻe��R$�)a�5~lߚI�m8�}l/������(Εr{�T��4��A=����@ü���,3�2�x������z�-U#�h�~����)ݲ���t3��O���5?��?��;ɋ�L��Q{��Zmבּw=&R�`qup�����BcE�@n5����O���a9"ɶTY��O~ԣ��aQT��p����ގIY��A	��^� �E|'� �!���E�^PVQ>\ � �[�-�CG�I)��0��>�(JWv\�"�^;�����7�L�u�F|��ð%�1t;�&a#,��'
T�DhB�����[�M\H�D|�h��=�Ay�˗/3�,2��'�Rn���Ly�١8|,ʽ�>�a�/z.Ƚ��||{k�}���VB"t��pZ�Z�M��=�Ha	��1��=�я6���3���po����!��q�0�Yą[��LaK@n�;(x�0�LT�%���F��&��p���d�jN�jr�4$����u�=�L5���!m��=ؔ�oa�L���f�!l{b�8N�4�$���AVo<i�g*O�\�4"�=Ԓ%7O{����T�=�y��ع8{�Dsay���'�bQ�*�֐�й��`�P-���c.Qnʐ&�F�5�1N�ܸ%���p���Ύ��,��jwr�B�*���kK%#��?�b�����ʕG׸:a�.JJ ��ʘ���!�d}a�7+X��˂g�� �vI��[��E?���Φ��=�� Ԁv�O�=F�@L�V�3��'���|�q�ײ&n����h�}A�2��RM�_(f���ڥN"l��#xr���8%2X�B��g.�qi�z�8*��:���u/�mGa~����>ق��#!'VT��7���    IDAT9x���K������M1�I�-ymD��n�Kh�(5uOc[�ư��2���m� �ߺ�"̌��ȗ�x�)��I�]�4�ys���y_���X���o�fj�H��:�a�S��<U�J��B5��wZ��~�kچ�=�����&z�N�
�����;6J ]�ۨ�2�;�t��L�c��<�F[R
 ]��e2ʉ�q�$C ��;\T�E���M'��|�GD��	�=�b:r�m(,��e]��',
rZou��� I�~G�5��Ae<�O.,�)����Uiy�g�i�M�!���z����x^�t�#���QYF��KY�;eK�l#˒����1�������^�o�gZ޶��Y7ꃈ�+�D��0r_C����'-�3[�Sc-g��mc��V+���~[�4~�O�k..�=�I�0��;4���[���"�ڠLJ2Ȟƴ��\[�6Y�ʨ{Z�}�+�U�rƱg����l��.��ij��p��#�?���~[?��~<��'UV]�j�PR4a��8�#��^`���I+�tT#M[Xy��>R�M����L,�)�?
ז'��:d���:�n���5��ER��M����zDgD&�l��<�k	�����<�<{�9�=3) �#3���,C(�`ȑ��VW�B;�/��O�uO�����/C|� ��p|psn�c���m�ڣ,�xb��r'R��,b��%U��5:�*&��o&�ml���{f*�r�ȼBtt�Q{�eѨ+eS��kaUJ}�uһԡ�V��
��>11�[W�(����&y2�
�7�q�t� xAf�&�]�,��}<�@��}v� f�]:3������Y������v;���y}s�;2]�үg��L�{�m�4ٞ��������P������N
�������H��:���%ix�,GЍ�G��4�Bn�t�愸=A@�Y!&/#]�
�,t��<U]�Ұ}D��LKMy�%D� A�)�`'��"r����P蕣4'gV����PrM�#�m$J&F�S��S,��̜�@˳(d-�S�kL:�,�;��G�2�B�H�%{ߖ��c;|�V�b��u�*�)	釭\^�{S'�Kǌ�pTsN�,�|P7�dY�6ʄR��T�<\CSD�mh�&u���< �|9�`ƝF��sQ�(T��z��z����dq�T��{n�.�D���rQnY.�ua�j���Q��#|-�I<��H!�g�Q�oJ��Wu��"�aE�%\+������sS������N���9�do��̈�R�N����V���!�4�+����)ZS�E��{O�����sT���_RBJP!�g墦C��v�����Ѣ�Q~$�PxE}�ϲ���;�<�Bю+s ���X���u���:$(G �Ҵ�@9�{HQ<L�%��1�D�w���	�|M��`"����@�"�rq^��e"��\���$"7Α���)���Xp�����QӨ�$05�ƚ���1���n%���~�"��iҶ�GX;���+�&��:k��Y?�%8"��*{Gy�6��^h6��]���O?=�ۯ���"�˟c!7WS�[2�}@���B�Jz�����i���-i�pk�@Y�LC�E�mz��9�m�p�#�;��3�2��aC^JN��#P����q�O��T�CJ��#� E�!�pw̔��"|�˚+E���Do󑅂eb�9MS��Š���14+�Sƾɉ��}�Z���a�-,*�R4�I~����P�KU�ԓQ�i��M8����|�Evق�U�H!���u5Cm����u+�y�W��(VJ?렟�6C�u7_�P�S`/2�	,��p�V�&*����oR����c!��佽3#s���Cd�H=)�����J�
�h�\|S��~�dX�h���ïMC�ՑHJ�[��I�����I!������*D�[�5�Q�g���[���>X��j:Ƭx���N�R��AS��o�u�����<�X�$�
,��P[Xm��.ۤ�C���=�x��
e�y���oE��Q*4+��z�����d�E(�4��U���İ�;I�����5$����k���MA�lӴ-�5��&�ֈ�Y6���
R��Z��6�z��s��!�
�;���f�>�÷�s,���Do�L)��܍��؈�3�JX1��0"��T*Qz�ˊf"�?M���$҄�m'b�p .�M&9�� P:w���X�	���
��~��D9�wNs�5Rs1�o���A�b�#�Px��{�_�?�%�6�L=��0ދfb���@H �H(�k<��� �;�И�2�r˺�aw�G�A�=�mD����g�=T�\��6�E.=���9�����l��fd픰d{i�)e��,�Ɖ�m/K"�Ѷ�0�/�/�Rw�g�0v<Ag��T�Q��{,�f�&fBU�C�������
[	�O��)�e�Yx���T�r�Y�"��fG |l�U�IF<�W�Q�/�����n��%��G�����>�;\h6o��ȵ�k�p�8�r������ԍ(��.T���^���ə�� ��l�l�=���-T_�,�tz��-=��хf����oI0�Y��E�ogvW;��ߜ�*�����68b:�s��&�ٯ�$���ɤR�Pz�Z�B�K�R��%�b"W�sK���l����7�.=r�(���"G����'Ȳ��v�A'���qwCQp� �Ny
���*�j�0�M�$<i�e�
���ò��o\%:��fݼpu};���3l=��'&f����[PL7��ds�C�~m�ե'��%�E��D��͆�,��] "P�l�b���qb����!l=	m�DD�:y�q6N�h�}�D�g�! ��t$@��b�v����<���GSD�w�#E٥��;�_�Z�؞L$��Id"�cg.X�1�(iy��:Y�tYv�DjY3B��<��wZ��'({8!3�[��H"��д���I'�(ID"�".�M���Em6�N�C�L��<M�a��,]y�E���tg����y}��Lr���&���E�BCxΨ}��X�mt��1i� Z\�����t�̙�K;��
P���2i�Dj�}Ԃ��	���`�]z�] �%��J��;1�q2�xC'�HFܛ(�(��e�<�[�3��w�|�!~�C�~:����O>�6��)��:�����!F�¦�.�
���"uA�9ڕ���Pg&�¬lE#qD��ә��\qRr��M�6����n-sG�s���s�����!?�B'$��0ѹ��"�,�ڞ�!��w��v���Q]	�#k��p-���k�k�vT;��Ȭ��[>��A4��{nl����׮\9�KA)5�B��ݭB"H�L	�����*�NlV��J�F�C���\R�(	?�����6���'��&�����
��^��<����g���yW�|��)��b��=�.�Ih3�����'mHW#�����b���3��ӡF<�RD��66�&(��'�D"~����וp�1���_9�av�֊F%M����G:R��d7�,����D#�(����i�u#%+JF�7g���tf��r�����Й���Ǣɏ޾��j�><�����b?�bY!�
g˒K�h+l�Dl��aie��ݶ��/r�#�������Q���eHdag���\��^j�OI���$�)YT �'��0�FK0�N!��"k~'⚉q}�$B���;�H/��˯��j�/|!�^�f2�Ss��z""�G�y��8�Ȩ�7���킐� �M�]���?�J��m�8��|�=�l^ �=p��86�Q�] +{IP9;��@O�-���䫿���HPxu��=PQ;��шJ.����5���t|�BD���tӌ̬c���G�	������$+bF�Ng++�a�pB�-[����ͼl�|t��iDn�4��[��,v.���(�q� �u�uaA��Cͱ(���l��V�B��,X*�y������N����H~[�D�H��"�)v���{F��k�Qh�YF9��s�8qT"�D��=���8S���)�G-Ȣ8y��/�{��.G>lnrq*[���\�.��c��J��a�INS�2q��TaH��,)�E=[���i@�bS^Ev¬P5�o%�iڐ"�1�4X�@���Q��d��zj�x���v:�2�Sd��F�&{�|9����qD�)�Sq XM9J�E2�v��ߦ+����iٹ,����� X�#�1�i�蚨#�n���`A�O�ώ}�k_�~����/�؈��9r �m34	4y��:����з-���!�F��H�F	�,���G?�߇Ø�@��.qè�\E��F��C�ú�����`�;��!;���skو�H���TEv����Z�6�o"i���5q��Uz{49�-.�4�(Ԛ�hv.Y�,AnǆB�ccBԫ��2��ǑN�y�ƵAE&^�.}���3��7�BI�O��Է���l�-f�4x�|.�p9ϑkȾ�޽��H��=:����w)��U�����m]�*�����m��A�����L��W4�Z�G��\{����k��&p�
16���3&�pO�~�������HN�ʕ��m�qXȾ_3V̂�XH��́��Ʊ!��&l_�#ņ���$C�p��B)ʕ}n�U��1N$���{��o����b����@!�^��}����1kc�l5c�,{�ANr��JL���z�c�b��%j�/4�����f8Ԓ2�J������FƳj�B�H�Y��]��$L���1��s����G�>K�
���z*��鹛H���<W}�ki�4W N�u�� }��Oe���HZ:UA#�t��<􏼈��mj�ac�t�.�~�&�J��8��QAB6�t��X�vwƾ��o_{��gK�tJ��=��	%����H�I�("ҩv6@ܸ6��2��*�"�5e�K�eŭP��$$Pt�I`�@Я �,�Hnh��v2�ϩ�7v�8ӈ��I�&�^i_�-,�,���'�4 �8ԛ=+���Nܰ���}+w�B�9��MlZ�ĭ
�̞k��c�">���1Z��f��Q�3:��1�$���]�h�.�s	_v�f���A���������߈''�&ᒰLb��l,#*��!,HR�Clr��:��:�
�r*�$lBBc�$[MR����]:�~u��w"r��m��d��w�X��zd݈�P�r� ��i^|����e"�},����l�&�J;�e�c52(ew�I���(��C��^j%�����wm+h:�.)+/�O�>��������i�uD�8c�qG�2�i��V9Ijǭe�"�T�]7Й�à�H��~�2W�^�֫�+n���[͐Rx{Y�l 'i8�m��'E�Y�a2��\���r�dNM{(=��)W������hٰeg��ԒNva�@#�[tB�E"M�D��C���Dh�3��hvd�<�b�;�]���]���e�ܾ�1�ʴ�Q) �?��K��!J���Y�L!����>�^MЖ�E�1M��%cD�n~H"%��K;4ǃ��]�EE�ߣ�Bo������=tg���St;�	�O��a&�J)I�`��/�3L �t��MW��'N�!��NL�q���DC�����p<YR��R�O�3�<y�@WDA\O�b��YĹ��A�Y��G��0�EZn\%z���	��q݌}���nP&�n��$'���<.��&ؘ֗���7���"���z�O���D|��'q�c8�-���xxO�݄(-��L��/\x�y��M�\o�{�&j�����{�`�m��n��m��eЮ��}X��K;�(�En����A����#w��<eD�Y� �������;*���4ul,��;�X�A�K��0�Ҕ�.}QwG��eNw� ;�=۳-�ω�îq��.���#����e{�r�� ��噳*�
���']&�JI�һh�)�i�YF���f%����t��L4; ��Z�8Go��������'�Cq���5;�z�7n�'�ބ䅎�un�ȭi��'l,O"xڲ5�s��"����4�#��D��
���0v��\��{7��Kw���*,���e�q�0���'�k��Þ ��&�L�RG����x�u�4Taʸ��-��>��yj0����ԩ� Pgd�ۍ�!�7�m(vQe'�T������~�#X�'�7���=�
q�e�k�{����/��x��AMX:?Ź�#�Om;�����C���A�\͖b�@�ゎ�x��=�_��1��v� Gc�$��l<�i~���܅'(�"��,��:/����K���-�t�����x��=q���S&�Ym�ʼ�Z٨B�^�����%�;B*ϟ[�0L�)�I8G	�Du�٠�S�����^��d,�V�zu;�%����01��k2ϴñuO�l����گ����:F����D���Q��L䎚u�RJ{�l	KڻF�
%:&E ��<�vR{�`��J�{�\)�yd��|� )��a=I��ׯ4��+���]?^��ȎA@�)�HƩ���)��EV�r�U�ˣ�CΞI/��\"�N����&��ҁ&Q�:s�C�Ň���с�&�=��N$�l�)vQ���E��J^�'4�lA4OA�A��)7T^�[&a��	�ω�:��c���(��-�ě�B��,�E���\��u�'$�� [�������g^i�-퀗0�ɶO��6n��t�}d7�ac1�bw��q�;x3�I6��8�b����]A�qVJ[	J
�u��v�����k���PC�-��I� ���Y�ҟ�<�@B�1����R����Ypmݥ{;�35<�7���!������-4.
���3�ܭh�[(qp�����in�@j����̙����G`�. w_�p� +�Fބ�g���2���(����I�`��A���T<�]Qc�t��X:�pK�y��bP����^$B�c�v	�����F��]n_���_��n��}��y x�N"�j�R�x"��O�_�e�=Cg��f'K������c����ܑ~\�&m-E����s����-�$)G�:(�JRq�e��J���iO��)Tի �ƛGX����w�0�,�m��Lە��).P]8��p]V�:�x�'TV]HPT�[9��m�R�2V�����P�Y�!��ԥ��(
�&O%"'O�cO�9�=�*��8cP�R�LP�<e=�-�,��D����}�(,���r����tA*�^Rm�6�x�RH��޽׼��͝H
�w�n܄y�$�>�A��m�aO��a����������.>h8oA����?_�#\��I�~��]�)	��v}ksdyee������Teu�P�(��K��Ah�}46RK7ߣ��y(d��� �&���8�`���mv�Lr6����_������]n��l<��T�q���͛���d�`d�f������tX�������[Pl:��_"o��ӳ=F)eA%�;exa^����Ű��&�1�.TX�ؠ~ݓ�#�|�قUP<)E|��b5��"6��c���;�����)�}K^�f�{t:�J�I"�]��L����Q^/�݁wF¨֓�B3Ǆw�^�YB�}u��3�'������j����f��]ξ��|ؤ�uGsWR!q���V	ҳc���ĄR���m#;�����M*�-��ǚ ���$qº�
�F��]gpn��؍C;GtR�2v�*m<��s�G!x!��,?ίk�jlI%��HNv��;\��Br!�<c�t"�
8���������,�GOn���#Peq\�`$�b�,�믿qՋ�ۋWmt����F�q"�`�2Q,�KB%�xS��MeH�]��>��ʈd�m��2߀L��	��z$�g���P��`Kȇş�i���k6�>�0U4*/^z����ԅ���$���M�Oa�#�nN�U�U��řy&���o4�\����*��YD�w�%Qua����#pP�L��[�m�O�Y�����Ѳ�h�]��Y��!���A�p����KKG����{S����B`��    IDAT�$�KGd������� iGl)|] ��c�
H	|��ss�{ڋ�/��x�D�_��_������.*�d�J!�E��. M@��¨�Ã3Jhԩ�(O�4j�ʜE�I�SF(ҁ�y$6�u��MeP]W,��u�c���;�*��T�{.�w��~�]VI�2�\�'�������c���/a�щ�HB�o��Ǚ#x?���o0Y���5&�WB�	�\���U���f�%�+�/�=w�0�6?z�Zȷ)�2xt�3�z8�Ԙ�ؖYN�k�ᵋt���i�����^U���K��X��mf a���~�ڸ�u\�4``�B,���j�-D|s薌p�[��X�/�`V�(c%2�av_ �G���=V�8�5FDzN�T�w'��?�����w�kv�{f�;�����j�y�y���p>���#���Aᧃ���X.��eTD��E��9�:�DӲ�	G*R���L�Ι�͛Lޖ�X���\� �,�;y����-���D�&�gf��F�;��Ǝ ��oG����`�� ��Ӽ�Y�?9E����l��A�䓟D���%�_e��F���7�T-�Ă"�\X ��>�}
���6�#�!a��#�B�4�s|GmۮB�0"�D'��0Ϸ	G��~��ܴ��5q�QU�h���&}�4+P�6~��)�Kl���cnӊk�SJ3�>G�B��<��1�a;\�@)^��������ɕ�g�]'��<���U�Qv���>Ԝ9��L�\���\�/�
��O���ocJ��NT�2Q%Uu=�oģ��0�.���B�sP�׹���������O��^��\찂��ajj͌N�����4~�<H�d=�s�	�g��v��T�مMR�Gge�͛��ߺ�d���4�$��J���?h��G�1��8���9��e!�Z+C�*mi����|k�//m�t+��7R$�q��?������o�.8�/e�VHv��cϑ���D�,[jB���c\���%B��d���x27�k�f��@.K��жW;�y-������i~��~�;�_�F2.����c�8>OX����_Dķ@����uU��+W���pr�@�=2!&x ��M&a�DXEaqc����[R7=���
��[�IK�7��P��]��Fѻ0wU�E�>�"�P"���Lx������7����Idf�`�k��me���{���Ds��Ǜ��1���kq�<�� )a��JJ
Ֆ ��ؔ��K9�� ۰V)��>Q��i��5�6팧mZOM9�)�	G�|��#����[b�Ka��Β;$�q��s�@��_p�B� ��{g��mT��M��{~g��qU�+����"������ٵ楗^j~�7�9w�Ls�!.��e���1nM�������;�_�P=�F�RZ�xd5,�`Аi%�H(4[n%��Mfb�t�^w�Fy���<+�"G٦������~��A�
�)��Ov��ń�Clʎ�e�*�y�8j�ۨ��F��L����N��Lrw�?���/�Q�v� R-?��&\:�.+��>~�[�fQ���&�}�_�m���o�u"�A܌8�q���ֱ<�!���:�z��݃	�fe���P��]3��&'���4�;��Z%�.�l�"6L�@+���wT���A4������L/Ø��%j�EKJ�a<"�IPT`��r�+��߇R�5���_r�I��	��h�$o�����3)c���U�&���1�EU`OHoTv$VT��fcɗ`h�c]���t6�Nq?��m�+�"����l�F�P�����@4	��&�O��&��0y82��8����VHE��/�ʪ"�JY;,
ua�6`Un����\���B�����b����pM�� ��
O��]��=<�����Pږ����f9��y��h�{~k�)^:E�I��c���	�԰@��v�:7n���d�A�H���~���&=I�����8�>����]l[�p߭�ᇉ��O�$����ߙ�n~g�	�T��!����`=���{B�f�/}�K͟�髰j��j�)U��b2'g��E�O@��X��V=��F�BƮ��j��	\?�LZ	MR�,\��Rz�AK�aQ�U�M��<5	����`���e���K����U�"<)���"���Jʍ���F�A��ڈ.
��	b7��[P�;ȹ��X��<�ؓ�����n�дܼ����F�
�Zmm��� �D���529G���}�d��G����i��G�u�oG ����D�b�fg�����d���@�d��1K�9&r� ������������.�.��̹��FE�� ���țk+淶F7�A3y4|hڠjT�4LY5���7�˿��(W�����g���t����ʟ� +�� �L�<|Q5^���_݈[��;HdV��
H���-/��Eˤa)�TG��Ƒ��|�In9������l���7b:��Ѫ�IY5���z8�U�ue�mpP���EF��\~�-p�nq
6�c�g����;��c�V�3�����_�~����(Hm4H);��'�ز¹�D��k�wS�]A�ҾuZ�ƒߓ�����]��ī �`�u�ub���JKd��=�2��p����u���\�cs�R�_k(P +׆����{��V�F���� 09�G��t�xh���e؈����q����o~���_�c�qq���A�6�5��Ų��<H�0�OOAڛ�ڍ��[�����#x|�e��j<�R��Ҁ��ičmf��`a|��C7�}�^C���
�È`���;2�k]5U�:g��|5�{}{y�O-��1a܃�n�������赟z�y��w`5�X}
9�è�.ѡO4_��>�#'P�� P��p/D����6(���G�z�"ڔ6���9e9��}W�Y����9=kosks���}�2��㗸$`�8�%P��ytss�� bS�ZꣿҔ셆kcE�����n	\��~~��"���X���{U��p����}���_�|�7���)9YXx�	ʇi|ON�>�ô
O(I��w�����a��My|���nj�Έ&6#L�%-� ��XDY��I��$��۰8�;e6�RﭱU�<�sU��]V��p��?�����)�ҟ��K �n���W�h���(�#
꽷;�|��Vs�:;�鬷����0�H-�(C�L$��a$�~;���Zu�8ܯ���>����u��w���V�?k94��\�u�Wp�a� �$��Z�aw������@�IdvWNj6�2��q����E�'��}�0x���e��;� $V�l*]�����H�����?��PM� ��qg��d�ć~��~���!R��<q�,�������н�v�[��"��ܥs���{��Ï����u2����*���65.�c0+G#���]v��`������b��#�A�)ܗ��������1���*���͇/?�&���{|@�6�������_i�M<dg��*K�^E��k ��bC�������_T�H?���@��S3��`���#{��b�)��bn���'�ߎ6�B��N��}�

�Td�dr����Ϊ�bA���N�$�fq��>��ne�����]��w;�(opЄ�8��dr't+
ߏj*���_dQ�f�}_��N����� ?��U��\���w�� ��`'�x�ѧX�9�,]{�Y�}��F��&���ȱQq���1�Un����ܜ��q8.u�S�.L6Y�f�m�5T����w���Q��gP�E�wuce��>���s�.�����h�\};��MM�h�z��t�x�u.oz����E���-$��� f�	�	F4��XŶRN���BJrGP��:�ui;B�ǲ�}K�O�-�<��p�� �%r,�fUdg��%E�� ��K��Or�Eg��lЁ_ܱ���4$�b�'����ɳ�8����������'������PA5�6]P�<�-W�e�(�տ�����w����/5�=�0���i�ns
����mx��P4z�����x�y��[L��u^e,tY������1�%^+�=�W�7�X��;l:VG%�Oa�I�=v����0����܅�,6�o�.6�Hw��B�ݵ��ņ�吜\x��'>
�\�	�[o��|��y��7U�3��H3Ok�+�!�Y��	:�@��p/~���1�*��'%��g4u���Qzc��%�(�lR\�
p?��?�^"9���J&��9r��{���(�OT�V�����h�5\�؉��/G!i\������X���=��6-����d'�A�<� g�"�mo߅M��6_��d��s��<G|��;�������g�����#X�h�����Ϟ�r�zIg���de�ns�]�O��7@�7��;�P��d�9F�	*T� ��1�i�w]�$�ͥ�97C�a�f�+9w��w�xͷ�����?D�{͕7ߎ=�&��kO>�qTw/4/��F�ЅǛW�����I��+�Ҳ�~�|=<�r}�Q��)��`K9��#_~�ؾd;�T]�#L��]ڿ�uf����4�`��fgΞ�=����.g?MЦ�|�9r?�4�>{ʔ�r���w��M-.���5d60̹��@H%X���-�9!Y!�!�����l�@
�O +M�H�d&Y2�/��oTH�Ѹ^�� Sf
+wʩuwO�;��c�������=�9X���z���Dl������c�lC�<�j��z�I����:�\8�p����W�ջh"��iF��<��{������wY�tTpb�̺�=Z�/�5��l�~�4�ف�G{ԳXPt��t0WYY���=���.����WG�kWO5������o�f����,�~�
�o(���@�. ���77?�Uý $��^�a�?$D �b�D��D�tp�hwޝ_y
�ߎl\&�d>�5�c�j�g� I $�ۨ&�)b����7����{I)M��x��V����\����&:�s{4Ю<�%���m��V&�0i ~�ʂǕ����6�t�_�q3��ɰ���>�	.rV��?��4�=�W���K��|��A�����2=�Hl�Z9�\{�G4�Xs��
�p$,�<���m؞E�X[]n�.�
x���N�+�q沼ƍ��|���7���4gΝG���h+�6�Ї�����eGJan/�B � �S�6��� �������lmQP'���f��׿l���s�E.���ĳ��pI�.�sT��m�|�8	�L?ä{Q�*�St\m��nJ���J�s'WkQ?�L�������W���.�n2ď/p@z��)SS,:LN��ϡ9%O�C���M"}��]V�B�ܥ�S�a|���3\�kk2��U~=fN�Ņ�(E����}&�������泟�����[�6���	��� B�Bvj�Cl1Xm3�{�Ή�g��<DgagM{k��?�ݥ�VA�E�G=�������-������2�b�����?K�@T��ۻ�2R������M�o�m�z���^|�N�$|g1-/�Lpq��$��� ܄}��>��/M�g{����SX�fy�V�r����������j;S�̇��Cn�m��$���ڙRc�Q�;3;��qoy�mH{���P�"J��-;���
kk�})nx�?�!0�5	�3�y�{��N3Ͻ�o����ΩT�|���_��|��h��ȇ����O7���������Os��$�>�\��@Yذ�����^J���i�Y�c�P>�L�yy�F�V��MOrM�z�4����+�4��WP-8*V�����I�H��~��0��0�$��M�����	�LL��L� M���s��?�J#,}�,�g�����v��~�6�)�Q��q�¶�2�r�5��M a",AP`�9.rCb�ҫ�ؘ�;�x�^�Ն��1�Z8{f������f�+����6�D쌛��1�_�|�P�W�JI�ƺ��L��.�a�������4���������qs�҅��?�)K���9��N�U$rh�`�ץܻw
����4y��[ל�r�H��]N�e�:��Y��v�F �H�2���N�
+��v��Ύ�A�]8h����2�:�5+�N>��]�Mt��k F
>��m�ap,��F�!�2-C�6)�QM?�p!}�e��H���i	=d�ҥG��}�QD���흲s�M{�ul�_o�_191��<���� A����̘4� >��w��l��-v������2\>�'���M㷏��^�2Uܨ��h�IIfX�t���o~�y���a�d������ͧ?����s��󋁬��PTTHY�]�\ZZC6~�d%�R_ܫ��6��}�.�Ŏ�]&M��W~�n�[��`����}c�C�ud�xY4 Pz(7T�r�	�&e>1w��X��Rt�K�K��#2	����^?��>*�:~�6�)Į�E�I�f<���x�s�ɺ��31={��D���<G�92�������U�d�����I��S)T#T@�Cӈ<��A�d�ׯ��V���'3��+�wӁ+�)�&g�y
�j:�lp2�z(�Ȯ��4����Ss��cPՉ���χ}
��S��4��	w�Oq}��a
EG�>ù��(Tv����x�����U��'Sy��w86&W�pQf�� /�Q9�.&Ċ��g��U�wx�������J���~�[ï~؄e�ǧN+"�?鞶Ά�W/ܤ���izq��Wp��yn9U��ܹ�9������b*�S���A��>��>׹�q �4���B9,��M
��OX)ˎ�
��+j��7�_׿Fd�u��w;���w��v���w)�[X�B��( -+�S�ҽ���
��ߏt_��o5��՟�H���w�g>��泟�,�"�:�3���Yi���&[����f����W��|�w�������C�/����,�c� ����Z�(<=|S�*��Dd7@��(����t� �����O�j��0�:��{�lZ�@{'��.Q9�C;稫��ťK�Z��^\.�R����{���݄���Z��|���)y�0bDj��bں�॒�gE#2?����2X�L?Ӎ��`��1�o��d���H�^P.�
�
�p���&��F�ӥ�<���[���4����������'>��,��YF;�g>�S�3�<K�x�����k_��P޵���p�ɝ8�vV#��V	,�n��K��� G(l!
�,�0RN+�Y.\�D�:֡�]� �m�$���%,¡�1��I?��w��3h1D�tK;��Vit���'�^g0]�HHYB���+W��?����DH���ٳ�2qF�ћ���Qj2G)�{�":�QunX�`"�&��w+#`45b�4��J��0;;�2���"�j��>�hZ+�#Vq�8�q^TF7�za��P���7/8d��׿��X�Yo��E���v���㗛ˏ^n�g	������
[�)P��p��R�3N�P���ɲ���s����������,�c8��E���0�+	ۂ8	'�M�׶���d��=��^{f܄��i"n�Q�)�u$��]�rz�W_�
���G�>Og~d��g�,�}��mB����ۂ!�Ʌ����d�V�D�t��w��&�j���>*|ݡ�8��v�x�m�2��|A��9��*Z�=K���臨5(��G����m�[yEny��^�Ҽ���܉�mΜ?�$U\(�����Y@vl��"g8��e4q� H�+�v݀  CX��C��nvʣL�$��c���w:�a�m�LC7��N�-�
��\�ZI��E��)쫣��L��`#'9�i�d��y�[����#h"���	#8��+�ʊ[�xĖ�|u�֩��;�?,�����LC ��}6҉L�����GbšR�bX���(��qM ��8i�	��Op���8���ltU8c�EG��Nz�	l��RA8+Tٽ�^��DHzY�0�-.u�N:��}3#��*a�߃��}�[�0iZ�������U�C�t��,|8=8��I���7y����
��Xj    IDAT�:.rC��!��C��ua�<.l	��iL�l��.*��U�^p�B�
F�~�>�³�1�^�wV?���~g�Ek%�_�'"_4�X�{���@R'��}��db���pl�"��;&��q�]5"�\��u�#L���HGpC1
X����7.�
��^��Rs����:f�e����0i[�2��%��ݫW	܃��5��6�n�+��V��K�d��θ¦�R��#�mK�A��$�i�C� &L�Z�>#����p ��r���e�_Z��q'���,�O11����դ�~'Y�L�p����a2��K�N�4�b�( :ÔR�/�&�ƙf�a����zxfHH[h/QRB"ew���8X'yIw��c��v �)cn����@L���|!x����zdӱ�=H4"𐟄U��U=KZ������8��{������m0|���OyO�����:��YC�(lXa�ĻKK��X�����m�Y߇�t=hjd�̘?tG��B�;�V�P��+gE|��چդ]��n�դ��2̠����"r�qZ^/´iG�d��3��8�Ӷ���r�w�KU���bCG�n��N��@:Oܘf�uo�.;}�b�JU���z��/U3n*[��-���p%���/���Z�R���r/a�	��Z��l}[�6!�K	�o#��E��N�p�'��K�|L[�W춠VO	�+��w������\Qs�(��.K��ذ!f��V�E�F���%Y|qX��hYP��6�7�a
P�=\��%��|�a2��g:�G����gZ�1J)�u:���"��Y��$k�.�L�,���cޠ��W����S3!
J����%��ɥLN"�
ȷg�n�u��qe�UZ�;ʄ-�ηv�#��"eY�`�i��0�m�.�|��p����o�k�:�~���)�Jx���/$JIHsq���YAv�mcc:�A�G�cSnϻu��������&�����451���'�/*�A(��ul
$0(��PƢ��2'���|�V����@�q(�Mi���+v3��K#c���zR�?��F �Di�2qb,�%,�hU����gWM�K#N���$p����6�Cs��V�o�X�|�쑮a=�d{��c��)BZi����nl�(�W�X�,��9ҳ�i�U1E�,ݵ~a�¡n��>��������x���i��j�Љ�CX;e(�a���w���1=JCMAw>M��nolq��̱��tjԳ�'Bϖc�(����F �S�@2�QS��w��mc x������N�&��wڙ�a��n������_4�bf��W�C؈~OvA�;�+n}� ��2�V�!���8Y ��WsX�[���{�����"��=�h� G~a�d	�`_vİ��3L:SS��A�4�Fn�p��THr"E�%��B`G�̂E#�ȝ2���)��d\W�2��h��
f8��d���4Z��_���S��0�vD�#~I�_;]�y�߃�&�I��q3~���Ҏ|�G�3��3�0{0̃����a��a�s;,��T��)ÉK>���th���0W��\܎�����ds�kJ�1Εsa������-��o�bJ����m��gE#L�,?ϯa���-���`�t7\R��C�7��|��|�ߴ2�v�+ǍΏ�TJ���Y��˸��a���ؑ/�uzu��t"l[��~���y���3���,u��1g9�Hʹ����Zx�)�	b
I<��(g��-�A�5
!{�U:Q����<r,R�g\y0wD{!E��b�nAM�':��}Lô�����dڵ_����+o�1�=���e`/�.�}�_;ޱy�?U��I��G����w'�>��dxG�ވז%��re�>��5�V~k[�(W�Ϡ_�^�G���c�sX��O^�z�K�ޟF=Ac���؅��xo�H��sQn(2eQ���H4���,MaDz*&X8+0ht��{��q�����}0��oÛ���y��i���)��4�3�;�]��Mr3ﶺ�/!�M��@z�Nh�ǰi���m��&���@^��鵟u�poӬ�3f�i�skz���m9ĝR��#d�8�3���IC��d����`��F#	!�\��D4�J$�(o)��}Ƨ6	�t�oä��T��]��p�M��W���ƩM�g����O|ݣ��ѱ*+~�1��">M�a�4�rK��Ԅ݂*.�N��D�M/�p�c��&�yT�{/^ێ��`�m��dX���Bm���������U�:�������R;+m
���0�?j�X!nO��������V4"�c�d�t��:��+ Ȱ.����3=,^ϿM �h�_��[R�K�q2�an��i�e���|������r�wڃ駻v�e�xo�2�`ܬg�>�n\�"L5�.��i)#��/��a��3N@z�96r���Ǣ�x�E6'��<��@�XU��DP����~�DA~;*���L ��v��F�����8�[8���.W��?)��d����[��������=E��k2-��t2l	���ю���6l��μ|7M�i����H�jS���W�k�`;���	C�3����7�u���Pf��u6b��Bܨ�Ɏ$�E�6h0�D`�3zk�Α�ɱ���Z��d�0���^��*JV
ju�����6��ig������8�l��x����ey��'��8�n�緋I�ᣛ͒i��g�h�ϴ�i�y�P�o���"�j;:�v��v�=����["n�Y��2����z�q��u|���[�6�)�	��M00Cb3+���=T'�����N�<�=v�CՏ0�Gnd�/���߂�߇/�&��Ii%!Y�ao��E�(!��[�S ���n���vX��������m�:y�,q�7��Q϶>�!�V��G�L���ȡ�O�ɲ�����g���̑��0!�m=3�LCgœ���x����#���p3n�+�Kăm���%k] �*��x3�^S�u9��t��tmm>�:��C����S�m6Sx+�����(lr�0�%�U�1o�5�"��
����u��/ݵ�=�]���j��{����RQ�u����ښt�w�3���:��w�ӽ�o�����^��'�M/��O�yf�����u�7�|�N�m�i��(�rd�FNU�6�+�=tq��6Ϟ�~�#�q)w+*��A4�%���}��w':N�qA�
ʬLZ1N>�1�,�d��n/�M8��˰=C���U$�&BԈ��ie�3�(i�� O�Lw���5��l1�n#�f�C�^�(s[�3~/,�,�w�[��T�[�"�-�3=��h�w	Q(k�kg���������8��'�i����m�k��N(/~H�U�bB7"�t��7��4���q&�Aa�}�2ԋ#M�GTlaő�n(�P�ر`�Q�'Y���jx�d�0����⦿����rS#���>���du����W��nRk����n��ս~L_�|�4w�=�r�������]{X�_��^�y̝+�Pn��gR�N���v���s�9�s����#��=���e��;r���	���+G~ æ�f ��F����XAW��I��6U�tO��	�L��}ϼ|�͠{��v��3�nX��c��kZ1�gtfq��T����!������,S�����]�A�����el#�n'K��9�N;�{X�u:�_/�/;v6��t�n.E���)��Z�a�����%�%��1)2�dit���g?Op������4CI�m�*�8��^������~[���w�����n��B�=�nz�QS���aܡm|�=m� A�D�*�q#m��zؐ�K~۠��Hl�@��{�a�,�@�(S����t˴�=��'��;ߵ{���Q�v��а<���a<H�F���*�r��ylO��mV�8�]��sw	�}Az8U��fشН>1�.Az?��8;R¤\�F.�4�
r*��JU�|VT$pE�NP�u����>����'�� �1��Nʘ��]SO�q��$�k6@�x��)���5�9=�ʼ���!���E`��{���*�:nl<���ٔ��:.ZT����������Y�D��8�e}�q��x�<��?Îia舔��w�a����$d�ݢ,�u�����7M��<��١i�� N��%:��B���i<`����'h��7�=����Fan�X_��;�#ڡ?ǥ�d4���w#�����y��1�q�ݲ�-�S����l����4����9�V�o���Ŗ�%�& 3��O�5��w�hIy3��3͌���4�6N��{q9�7��=�Ю��u��ޝؓX-�o��'�_��Ʃ�qZ��H?3���薝#����V�a<W~��_Q��(ܸ���N('�����t�N��b��"��a����{�8�{�S�F�KhA����I8��Ev��V��xÌ@�q̓��o�H�6o�R?���.K棝�Y�9���43�i&�3ݴ���~��ߠ{~C�	�G��#�,�0JS�+��EpM�����0-��s�Gj��3^�=N:�kAG;0�ā<Q6���3��;9=���w�}��S��|��V "�� �[3�!a��&������=��m�fƍ~2,M����_����c�A�_�0� �]����������In��v�{ �&IE�!ːiG���"�2��Rg���F?��=~�i�g�%^v�2�::�t�]��f�דw��ά7�d���~���+k������][�`�r�
��vc�o�9�D�sߢr-2��� �"���	��0 Lҽg�n�H�8��A^��@hKy�o�밙W��w������e����g1�F��i��|ҭ�3N��N7�x�D�˷<�O~����_���y>�������6M���m�>�hX�ͭe�/��R ���o��,��[5�繁��}"�!�a��S1�vff�7]*uq��*��V��d#sT�%bg�Q�ġ�Z�N�!,)H�|�6���'#µ�v���u��}��/�&�t��L3˞��u9�{�?��|�Idlᓰ�8i��.(oG��;M/�<ZO��oq����.���"��t=�L�!0�_|q�2j���p~��'NMNL�ܾ?;7�[�A����d��
���nT����:=8�6D��T'�O;����d����ie�f�t��A;��ݰƷ��������fx�A��6����f�,����a�.�;^��K'GH�5�uI��-¶R��iK�J��S�=˯�q4q��˗C�D7ÑO��g��g�ǀ96�^���8�iT��R�%��cۛ["����H�X�@��2�X�u�1#�f>R��v�eH�gڲZ�r7��mD�!?uX���7�,������6����t>P���ii�̇�9�\ƣ0QE��巔9��FTe5�4�OR{�VD��tK_Ǎ� :Ú�&Jӳ��#��Dt�9>~j����G"���Q�C~�d����P.U�����o�MLm�r��9o��P&�������J��#'�D�
�[ �0��[��_6����&��6�,�ț�~k���A�<ـ~��1}��|�]��X����I���OiSZ�h�?P$}Y͂x�oy2/�����y������]9|�P���e\M���<(��+�&��c�l��p�X.ӊ�X�./�5n��.��E�%�w���������햍����?Ǧ�Ԉ] D�u��!d���qoทh
P�<�(��T�TZ���U�����W��_do�p H��i�/.}�g�mxJ�Ko0��ʐ����D�U�ֽ ���".˘��K�gx�f�?ː߇��yfd;�>ᇝi�ݖU�����i�S8�c���e�8D��N۴ヷ�Ep��歟����2��>6r#��S���x;�<6��M]��Np^��)��)�`Q�f�WX����A���z���DP� ��� ��A�u<�3�t��=dh��8Y��/]�M��'h�$�@�#~]��;����01F
���t}w�2LFd�d��W��-S�7�M;�%d�]6_�S�H��x�W�Ɇ�ϥ������.:���C��3���].S,HvY��rF��P>"d�K�"J�SF��AjS*��u����T�4|䏏���`���2\�#�3d�V����2e���ƫ��ib�}|�?�@ϸ�^�#�z�F<M�1�D��3T?ƕM�چ�%��h�^
�-s8�g[��_��R�0?({>~˺��k��rmm�c�����t�9>rsF T�;�F<�w�߹z�����X������De������l�D^�&a�v�m���%l�Q�K�/K��6N	[�����)��?����K���o�W+�m�,g�d"^��6qL�������o�M�Y)��d*fݨQ
��&���@H���8-�5n�G;�Ԅ0�ގ<b]�׾ѐ��5�H���لrd�H�Ȟ,.������	q�%�I������C�IA2�k)�������ٵ����+U����0����zŲ�Q��!,�����u�`�H��P5������@���42�v�>��q3�ߙv�ND����&��IEu�"N�L�ș�l��_I��-�A֩��|hĤ��*D��vVM�e�O�b��}?Y�,?��I�L�T��J�,�0x�7�z;��u�v ��@s�֭��ӳ�o��Gzf�a6sHq3N��5�\��qj�\a�+�t3�Ҋ��T!:�3s+�4TVZ�6鮛<7�0ݾ����4�=����������l�3-��hg�}���M�s4����Y�^z�G
�C�*Z�!ad�|7X]'%#��w�*��k��r����\�(��3�n	�˗/�q��Ery�3g��fKN����Ǧ�c�{���b����o����Kw�./�z������fc��Ie���R�,�4� �Ү�{�~�[Z�}�L��f�A�H�u׿��<:�a4���s����w��-"��v���j��C�j:t\mөM~�~	K���#-`�H�q2������"��uGY?��-3�}v����g7ⷡ{~m���w��w)��0��p�a]�/��/4W��aܳi�VW���D��p���ͱ����nq�����?���~��G��_���%�,�xyǁ<����*^��a�he� &�cx�]_��%���W������ ��,Wc���P�D� : rn���I';D[ j\��Y3aB�,�s�D���R��f�.A��e4>�"D�eE��R,�\&��x��	�mo�f�dC�g���ˍg�����	�b*�
�4�4GX`��A �N<H������W�� ��n'�p>y����(�G^�W
#T"s�>�O�@h������RG�R7�i�4��~�R�4^|p�扽��щ���0u!�w��X����]5����޽{���8��}�'yD+���������;��O`�i�/`5�x+���H�:G�Ѱ�N��+�Ӯ��M�	�wʑ�Y�ϲi;�v�n��Y�}�ʶ�?G6�2\)���l��)<{�>4v�o<�a�?�,_�~�a���a����=3L�~�V�~���0�G�gx�&KKKA�� ۸�4���M����#��ʠ\���3���\������A�&Y�^��ʻ����~�f�0+0�,,�!X�`�
��bC
i� $�Z���/��Eb�3�XzLO�L���-�rz��ߩzo���� �}����y�ɓ'O��Pu34x �L"TXQk�߻���5͎���#��ߒwL�$H�`�.�x�E����o���ʉ_���`9vފ��۬�DL4��X\�]&j���D�d�>��s�%����v���
8i�#��6u�q�Ӽ��p���ģb��Nެs�_p������|l�;n�e	K����i:����+�m�󷣻0�	�፧�k������T�{��M�� aS��c���}C���m�[�me�9P ���ޫA�u(�� H�)��'Ț Ͱ̿�m��qC|�9�n������ST*� �'�:�yQC*W���{`���89	��	��!�\ۜeґĖ�Ɏ�&���AÅi:�$R���    IDATz2�vQ/kk�P�(~\:��߆��EF�"��n�7�#n�O�7<g��oې��?�1L=wҏ��<�Qka�ߦ���7q�l/��>�&7+��ܡ���S�o�C�
�>*t+p*�%\��@Pb�w��!��iZ 9@ƿW�Z����P���x	e{�Y_�,�'��[F3���~�%�Pm�{��y9W�v.9�:)p�D9U����(�6!l�Q9�Sۦ�G�-�Z�KyN���j�j�B$EK��N�����Z]�1�i `���m�E>�Ƚu�%Hb�q�V�k���i�!�5�_8�����e�[{��o���0�ۦ�U�
�3�7J�M��76̌:n�����FG�6�  �#�f���qr�'; ɢlP4>=x�˯?�͸��K?�I���f���2,�R�5�tƱlo+ST�N6k��v�q�[˴_W�hsnwNE6]�Q��Xyӄ�Q��<�P��5�Z.0�3.��SG�����00�I�n�lk�}/�j�*�eX3��2M�3N3�f�2���WK;Ju�R�m�E�����qk,�s[s��V;�~�(Cx����Jg#�a�9u�����lp��Ώ�>R������Ęqrk	�щ����!u<�y�1�O��wn��Pc*��w�+����Ǫ�@�Ͻ��e�Cekr@��`��D��Y���e�9�%��!acT&�d�z3g�trx5V��~�3^�H���g�n<ȸ|�T���n>�4�t�6�ȷ7FJ~���c��Lo�$l;�D�O�6���v�p�%w���/����n�_�At�K W�����M�I��?ٰ��6<1��4��;�3�j�(_��n��������-����׶3��29Zpb��1�5�#՟���N�=Y�?i1.��].G*+����!���O<W_E�����r�b-�J@I�v���8I�����('�ǯ����r��\l'��Єg���g�a�m��M8�d�(�8�.����~�4��Ҁ���靃({[�b�߈pX�m�o����Y�ܖ�����?�t�؉ٹ�Yv1T1E�XyS��_]V�J�x	�l�a�峍���3N�D�@�pަI@gj�!�s6��oE���t�k���b>!�P��E�qɸ�7*�������~���/y�;ʙS'�[�r��yzv�����Y��@T�O����g~�_��7��a���M�P�,��n�G���h��o��!���O��0�j��/jh�;@���y�j�5o��EZe)]ԧ��߰�'���y���QRF�O�L���V��h]��-#ܶ�0?yة��[��[F��z�_&Q�}hKX��s�f�gʥK��&g&O��j �ȡ1>: �uM��8�g<��7�n�����_$|!NB�� T�@�1qR�0��.D8p�]������#,�,/�I6ʻ�����|gy�����F�=���A\�f�7р�H���n��ɢ�n��Un����������/�ŏ��ÃC���7ʇ>h�)�W�];Kg����m��Ω(C쀭�&<~���o�����4��m�$Ќ��ɷ����;4�q�i-#�}�Kt��Uƈ��Y��ǟ}7[aڬRm-R� 㤳����O�M���È�@�{��g����������S�P�Վ!�3>P�a�	����9���4���c�@ME���㮬,w&4-n�],�������a�������3g�F��;������t���Ъ%AL�Z/�+Kс�ۨ�P��n�@�̗>U�㻾���o����� � ���#߸G�vKW����au��m!Ǉ�����f��ſ�ᨶ������e�q�m$����5��6]0�x�N\>F�L:��q�dX�M�d��D,A�F���x�@_�@{re�3�xß}7�!��t�{p�Ņ��Y�=������К�͜��I'	 l��?�N���̣Ǹ��N��n4�yBt0�^�hSG�8-v�&�,©����ʷ������?/���x��ܭr��edt���=�텐�Gǆ�2HPk�ۏN{��^��^,m�#��gv~�0�5������|�,΁L��H9�O�˶�	�KOo�t���:�Ǫq���F�He%����� ���[M�"�R�O��~�8M��	� P��6��f�13��X��ۺ��������3o�c>�x�˚Ag㼑`�웸U2o��ͱ����S���.]�|�����@T�Q����h�g:��8��ЩJ@����j琯�6���R.5L��w�ÕZ�u�G?2v�d�!qjz�<:V~�����)O<�tp��7����H�mM�P�����Kޜ���\j)�ss�29�k
��7�5���|��`5�P)s� X���A��o� � ެC���.�;�sQ�
\��=���6���X�
�J�D�m����a�*�/�z���:�6c���-F��9�tF^)R���0��d;���\Gn�D�ށ�m�d�Y��o�6'
��,�щ���-��s�6�����Z'^YjT������26"]�gC�?߻�6�3����8	@�ã#\?����g�BY�+r�U�?�ߖ�]�QN�8VZ�}{�vi��0�0�K�V�a�ٰ�_(�䱶��|�P������ksL {�3��.R��/����\Y�X(0� |����2�\F��n�3���G)s+(f�DR.�dm�KN�K��n£����L�y���4��n�_~�G>7t��诬��E�)�����D�:<dO�o�V�`�����'�li�966�+[V ��a$��?6��0g����{�7��"O=q�n~��Ov�9�=9�0����|��{��<������-�mO<^nܺNf=eim��,VʁC�M$ N�,K�a�Ņ��K�(tn�[Y[(K���Y����UeN:bIԍ��2�����C�-��(�T�C�O=���V,��j�=5����U�Xu�f�颭�X%��7�%����;Z������:���¹�o]���|�=�UV�6���89�J�T���F����W��{n~�d�}:�p�9�z��Iy��-f�}KK�C�����:�A�Z�d6���iX9�9��Xc�L�O���ٔ��{�,O��K��dp�<8Q��뾮��/�<��G���g�0�v��,hJL;=WO�w��6���ѰeĔ����؊&+�p}k�q�hKBd�x^ڵ��qtx�\�~���^,��?�n�zQA�]�ss�,a
{���r���N�=S�H�� "Oߌm�vO�)`[�.`%<������?k"$�vǈ|:�)v4�J�%��iį.�,�wı}�/�ŏ�0vt��2=3]&����9��훸�v���n�i��GZ;42�422�b���BD %"�UW�X��y�٨�/|�;�6y�="�'�bz�6��.��:9�����ȷ�3�;�-���o��������������-?�3��,b�8��X� ��eF��!؇ö�K�=�\�|�}�K+�c7������Pk�](]}��@��� K�uu��i�Q�G0{EDi�_�n[e�`wz��8p�<��g�����K��G?�2wg	9��ϔ2��0~`��۩6�Y��.m��+�.,Y�#����n��� M�&bL����o�ո��$�:�1L���HO��h|7�PW9���O�f4#��#A�L�[�-�����RYX\ w�V���ӲN.O���M����H�nB4��f�jn߹Ӻ35}�ƍ��rC+r/�� ���fx�U ��o��Wxm�������p�$�*/ S_*�O"�_���]�*_�~��'�SSwB[6�X�4 �A\���OȡoܜD.$��M:�~�et��������#�aq�E�ۓUMj��6S�5F��h��p9��q./��[�7^���O�x����R����-�{���0�.�=r��KmW���.᫖�F��$NF��2��h3����w�%<+�Ubn��;␮7sI��̞B��S|����5?q�S���1D�eĿ���-\e`��훸=f���2����JЃ�]#�肆�v��o�Gm�@�����{��ߘV����,�I�����|L��&��u��ˋ��������Q~���Us3�����7�!�jiK$r
��B�=��$���opS�2��YB�1��-#��b��Vy�«�7��[7��;�b�I����cTa�����9D�6��V1f�A�(;�F��0������ղ�:�:�U��-�*O<�X�uy�������k�X�Dg6V��c����d����
c���C��ֶ�D�7�Bh�1���vʻD�N���1$�T,��U;��Tg��ša�j673#�p\X�Z��T��"���M�� �1�a��X�`p�P>0q`��x"=�F�ƭ��׎s�`<�Kx�W6�����ɶl��^�t���2���P)���G�G�?�����_�;0Y�2�0
�WK����y�g��z�.�0s��M��S�����r����g�`���j��A�GN+g>����zp�"2�P\��*Q�W��[�f�p���z���/�wXb"�B]��Ï���vy�3/R�Fy�˞(�=|��?���eq���m�
m�� #��=ȩNb-��C��X!:쿙K���?q��t�߻�3V3O񞋌���nA�Ue�$甌Eݧ����R|:�;{߉�eD��ܛ�n�T��׹.Qi+nQ�S�d��eG��"�w�P�m`d��x�c��)�����5�~�cE�w/�2� �����d��gx������?�? f�@��Qg�͋9�u4#/��b9u��;dr�&����1uy�u�Y+g�?!v����˅K��(�O.�xf3Z��c�)�G�����2�`z��5��AȜ�;`��i'<|�H9x� ��iĊR.�|s�Vy���Pa.�˯�/�#c����������}���⫗�X�̈́a���KBU&L��qx�/ A�w=����t�:V#�s�?�m>Y�6����iS���$�N��By��-DV�;W������ު�웸X�:�����/�e����X�7�l�oh��B�S�t�5N ���ݶ�̼���G�SV�!�"�f��o��o.?�/�r���a]q������/?V�#O<B��GE�9oay5�mD��r�ܩ�>��Ǣ�}h�z��2<1T�f�ʵ;�����L�0�Va� ��"dx8uϘ�౔�v3�숽ě`Yd����-�
��a���4��b���+/����+o��'ʍk7�s/|�|�S_�X�E���/�Ͻ�j�7��
QJbvBg/'ﺀ+p��Y���[�k��F'yg~7��<��bĕF����S�ڕ�exd ����o�N��܍�����}7�ބ��J9�;̳S���.��u'��w���-� 8��O�]�3��qI.���څ�P*`�_#8�.�a��y��5�������-?�S�c9}�L�]���/UKw�߄p�˷~�{���$\e	�y�ܞ�Ew�����O
���W�^-c��T-��*C��f�E!���xU�ܕ	%�a��D�b�Z�Ů������ˍ��W4��3���s��XC�^@C32�.~1g�0��r������k����˷�?*���(]��_��/ï�p��MD�U�(�rw7��*�T;\Z�U"6<ݽ1��ɰL~d��M��ծ��l嶱
�@Z#�7��p^�=�&j����o���m�u�:+g,��ғ&�*ہD\i�
�X�%�jl���w�w Jw2i��8��W>�������1;����So��������Ν�ஊ+��.O��_+�,��6cf��<R�_z�|�._��_ZN�=�n�r��Zƒ����X?�ݴ`gҶ$:�256*m���+�s[S����W/�R�#b<x�zpN�A�d	�����X�^�a�}��Ce��hy��G��+����}ٺ]y������WED]߂q�F���>������X��I�:j�n9z^	cGфa��w �?�I|���m��;�o<�����̟��(�7�k��˪��ʚUP���/��6��Z��)�"	����l��y��WƬ�ĩX���� ��-�͆[�Z������[c^�E~��t�ޙ�]�?�H�ٟ�9v�� b`>	\e�ThZ��uџB�mT|�Ja�ň�z�tY�/>�e
N��?��+�g�8P��h([� �8�4;U�f�Y�\@��}>;��b�s۶�v4�:t�@���̡j��Q�Ⅸ3\����1�tN��[��}��K��.^//��jy��g�[������gXI=T>��O2�`'s{��y{��-����t�G�#�쌎����a�)q��I?���[���u�|�g���M�>DA��<MWEv+������������=�~��{A�p���k�*6+�j��k���+�	���֤k� ��d�K���۷��%L B_.g��aLy�o9��YA��s?����w��!m>�˹�t�o#W�e=�E.���_(G���G�-��w��/}�Xyۃ��o��8�(I�a���e}���$
6F�~�w�GЉ�$ƦD�nԌ�c�Ľg��5�Zc.��?:!b�,FC���e|x<��r���#��&-/~����|�|�}e9���2s{�P�o��o*�G���~��R���PAv��w��a]q �	7��O���N�8#��:�}$d]�[G����b�:0`+Yı�۷�o΀���.B��7D�KU��d	�sL����B^db��r/�  ��p3��s�L�| f.����I`{ԣ����1쒧r�:6���� �����/��������{�ɐ[����L;��=qd���xp���-�k�A�}��b5t����d�B��;��q#G�չ����$�z
���t��Q�z�\���jR�Ս���[pDH$d��6an_��m���i������c|��Վ,-!����Ĵuji�ej�/�_R.�r���G?X�|����S��O~�S�U��Uϔ?��?�6C-�փz�Is���Ĩ�p��ĭ_f�?Zx�G[�h2N�#�#.�Y@��������[�$۲�TN"�A�>6::�r�F��Hq�?�&n6�`������O�b����L(?��c�r�>I�����!>�����@�u���L�o�3�^���Պ���0;�����?F�mv{��L,���E�$�~G��ߚ���x觗]���?�ɏ K��'Y49|�@�'��׮�ZΣ��B����h:�Zȥ=|G⎉2V���D�	�
��Tn�Q�:���T�F�t�W�C3`۴� �5��W!�j\�8x�H�9}��_%���G�'���v�|�g��o�j��+���[~�W~����kl��d`n��U�J�6��u�Z�^��vV����7���o��_~'�7��;�x��0�W�b��b�żzt��	�n��=҉�S[ �" +�۳�aL�P=���q	 �l���#˩u�'����_�k~�|���N����k�c�OS���,����Q����I�\�}��[AE�_dw���#e�=SfYJ�ӟ.g:G--f��3�0�2�tKM��0�V�vG�L�Xu�@�j�f�PB���E�=t2H��U]7D��5aD�m;�E]{����z���՛�ባ�ߔu}��By�'�j��+�˥[��S_�ty��"�L�Ǟz�L�b|����u]�đP�x:�Z�V���Q>J���:F<�4q�'d�w5N�%��ȗ��v$�q���/��'9�D���k�9������[\��o�^n�7U�"�޺y+��yn/^���>1b�3r�g������o��t���w'��oôs���lC��
_pRc���7?���=��&v�L`x�b������7��FO3+!_�6#����it���aӱ�A�,�}s�:K����Ct$�g�<
D�K���d$aS��"R�7ce>�!\�Y���4��h��1;��h�cP�ҋ͈�wX=�0���{ј�o���g�8Sg��	?�Fe�<�����#�ș���W^/��,�=��5�[�X�D���?��r��l��	�čL��u�W	N&�V\    IDAT�5�6�Q�.��m�fX����;eV%@�;g���˗#^�/ 3Eq��p�pwS�w������\�p��%+t�����/z{칷�I�6R���x�w?�0�����_~����0���-@��D��?�c��qrj2��89GP�V�я�fQ�E!h���?�C�Ҟr��1�Z(w�$��r��A�#,��D|9x�P醐{GF�h^*�;FG&�ɓg!^�*�:#�;���\�[�a�{��G/�^������},"m"֬l����$WRG �^��[,r��&Y�Y�.e��>��'��s.�u��W_cԂ����uy拟.GQ}R�O�Px�q�.��q�c�B?���;:�,��W��N���V9z�(�EN^��/qc�?�C'�7����7F���g?�kiq4ڞN���\���#nd��A�lN�+�;���4i�|"��������-Ӹ+��~��2t���V`q��I���Q��}��˷Xf�x����g�!��X��d�\�q�̈�bM���G@\l&�hx)�S���hvy�6jŀ���E	C��K�۶�"$�.Dq��X�uH�� ��01�\ԛ$��!������X�y�v�ڭ�V�5aPn1�@?~��!�$��#���Yn_��_U._�T.�!���&���o��7�g<ã=��t�#]�J|�<	%NƋ| F���T�:E�d����B,��ٴ��+3��YT���g����Z�*���u�!�Ǭv����r��;7[�[	eE	@B�Qx���r����$�rFc����� �+������ �mZj:�?��B��;W�����2���Y��W�m�%�vn"�ݙ�]&O`�U�7��?W��6�c_�X��Q���e��]6lI�c�^�w!E�E?n�\i��6:f�����Uİ�C�?N�<"^L")�{�:��l���8�~���:�?�mN��S���#�SNkh�^���EwD��0�]���<�m����O�-�?�jy��Ǣ/������>\.��>�N���d5���p�zhgM1�&����#���c�S�m��4pD���G�w>�|�I��㝂6�p�g�OcW�[}23���c/��!n�cо��/qo��3����N�!P*��v�>���h����x=4��S��߫nٻk�#�W��۞/ �ܷ��&�9����uo�6պ�)�����(7��pX΍����h�����by��M6,�DgfC��u�x8)5�6D�2�\f�c/m�u�����R��3�l	T� �b�Z�,��a�����26Z;>\
z��ʜ���H�7�!g֕M:���vC5g�l��WY���|ײ�0���s�4���S�~�Xz��'Y�����0;�PR��a4H�1� (���	{�xI�gr^�����q���㛯����3/�\��"©�y���,���X�][�A)jX�#G��[�o�k �����t���[�l��l`>��o�R���@nz����\y��u:���'d}��锹gf���6�Ͻ�\y�[L�yЉO�Yw�?y�:z�u����6�]H!Zx���7���Sw�%�E�ι<h%P�u#���mq��ۦ�׽�N�5�b�[[�艇, S��c)XB���g�0sa�sw���*���F���~�3&���7nÙQM>����/>W�����(���-o������ ���%�L���n�$>�đ��N���t7��wtWI��Y��������%p�7��f���/���]0D�n !8e!r\��>�����Y���A��葮H���a>�݁c��{w���4WN$�y��?��1�΂��� �E������ٍ��r��q|�\�v�vk5�-ƙΔnV��[;<kw-׆W��axU�F$�Sk�d��VUY��w��]C�-��~�#~��
c�oa3�}�ڑW�A�����!Z�9^ �l���̅!��FY]� 
},���"������?t��ȞNl�~�����ʱ#tX����a�_x�,#�n9v��:7J�'��x��,wkP2�n<ݝί꤁��q;]0�z3�LI7�0��`�V3i5�[r�}7̢zƞeo��67��>����Y�$���H��Vmf%���[@e�0��7"��c�ݡ��}�� l{���c�c�6G�D�Z�M�sp����E������W��Ȳ9m���n�m�8�V����О���
OèM�z�,t��J����Cs��݇ȱj$MV��w�j�$�i<�P�B;W���.�ۑ���@n���!p�U/��]QN��v!�r|c��W;����=p���U^�z�<p�2�>�.gΝ)/>�
p���.q�L�^��w��q�2xԏt�eG�%n�u(P��x��X
�v�&̛���8��� ��V����`�CSiD�&r��lx����-�i�f�ɰ�6���ÕFw��)�W�D]l����! 츽K��6.��v'�g�2l_G�
\}���D�]I7�,�s!(6 �Hp����.Z}��Y^nn�`�ǈ�[M���S��'�Jؚ�
�8�U��Yͅ�d��=�
�|�����ܱ1��~h;89�Ot���тY!*�W(YWG�뷯���0�������?�YT�'����?�hy���uz�2���`OHGb�9;p��(D�S���H�������0]�c�3m��N<��ϑ݉��u�rY|ۦ�f�o�:`x�Xo��"�8�G.)wH�0�h��٘l���>�	Wߦ_5ߑJ�G��f_���|��} T 	�:�\Ἶe8�;cf�/_�T>�z=��<�!��!��%���&���e&|څT��#R�c0"'��p�t�y�ܶ�Q��<�xp�?^F��YJg`�G�uT��>�B�tT5-��:�|�!��i�o~#�@ �w�ࢢ��v\.��C���6w��E�+}���qt����:o�j�l�]��h{��� #�b�6d&��th�r��"d��|�&���?���0��3�;o�+�G:��,l�.�<�;a�{�Ľ5>�օ9�G�HU�>{�lp	�J�VT��I���ݰ�w�4��yd���%}�;�*N\u3�gjP�����nZ�V7%�m��+7/ý��Q-(�o1�rgMplf��A���JH���q�25�A�ѷ�q^q!�4���=,ǐy��4��6Z�iF�ؒ_���"C��^B4�*�ؽ�́?����+������?�8���7&�pl��HΈC��I�ѻ1�y�P/։�L��f&cdz�	�G­xPmWc����8�@Bd
w;�m��4�M�\G��1މ?�~���<���w�'��`N7n�(ׯ_�<�0m����֤M�Nw3��~��Ĳ�:���6�G��_�5_"����a�����l@�ec}g\�(��g޾M�oӛ��l�yNc�t�/���"�+;4�EC��>ȉ��h\	�=ѻ"�%�"�ݦ��/bҪ�����D
�3�4xB}�\m27:R���A�X>zQ�ͳ���(ps�N������,�ϗe&zn4�]��7�Nx�\���\#��ɽa�n�v��x��v�∓N���qք+pp��8�l(�n��,@qM�.'��{��r,�,���@9�~MՈ�OpjzM2(�(�+L+!JĆ��čp3N�ķaMB׿�.���r|�0+N�\��o�kq�'��Mܾ�{dd����JX�C� pO���$D`���� �1�$N���o�y���Y9L�f�D�q�?:ĮA�'E�(nܐ���{Y�^�xV�!�qs�c)g�CE�ї�3�`O����zƙ��c��Ǆ2���ȔWm���pkb|{k�D��Ԋ�n\��o�;�e���[lfq�>��V*>m�
���/W��W���s�F���U���n�	�~��aeՑ�c.^�j?��N�+����g���2�<�����A
�g�w�@q3�/����@ša�G��4]������m{9q,�:u�T���{i�c��j���9����z�������+fu�*���0%��}��Qy�6�FAST�Y}�f+�8�q�O��?�w �]�r�U4��4��TF�)�&�r� L�9�A���������tp��FP+�R���P��^ۼ�������7V�'����y��B�j)���W��[#�qW���.a�@Ⱥn��J����AڸH��Ȋ�ת0t��o'���K��l��r/b�O����w�	��)�8���q���\�!�	&�m���<&�k�Kݿ#��*�����r��U��N<�����������y�o'�jJ\\�a�8����\�|o��K��?��	A���}c}��	E�V\�'����9[Q������&�鯘��cK����	�R���y��7~�7F\'fZ�b[��Y74x����Јx �;h���%u-����ۊ�W�U���2��gr�(rl�x |yq�+hK}�n���y�bF���ys.�*"��q���M�Uֹ;`$����?�g�8uJ�S�{#sR^���4|��4u�j�7��G���+�ۮ��Ƹ��fp�I��y�|���娊���8��5 a�?2���1G��y���y+׌�� P[���3N�Ź����:�S:��p6:�/��s{�#��A[��pP�w�F�ج�o��ț=׼m���trg��v��3�~�y�~?��?�&�r��T��c\ۆ�8D��]PT�c%���fPNh'��Ғ�1�+Vݳ8��"����������*>*�ɟ�I$P�Ze"��i�'��lr�D�N�ـ�	)k=�YU�M�u��Q�l�v�Q��<�r����HG�u���$J�u܍�h��q�͵'Y��V�v�q�Ѓln���	�g��=|XUj�E�N�n0��¾�$��'��ﬣ�L��淿���xQ�I��n��s���n��#�� en�ەH� �;w.& %V(�+���ƷWJ|>��Cg��w>~擝i����8Z�2�zw�(Y��Z�T�\5'KL��#�0��H�dzp��,�q&6��P!����I�N��&MZ���Z�8�n�Jc����R��M�/v��:r�\���p^�#��i��m_�Q�\]QMXȤ�A�U|����Ś��C9w2ML7�f�G�!����q��.�{�n�x����ʴ�ru�M\�N(�����,]�:����?��<�-�ģ8�F�W'N�W�YY9�'q�W,	��{�u~�=NK��iNG:�p��Hl���P��F�[i+o>w�7��Q:�����mfNN�F�4z�ɤN@̡�0m�Jױـ�(�NH�[���RX�!bH\N���ejy�^L���L�B�*���N��@�=e!;�!K����|X���à�3��Lԝ3�T����-�I$�@��� `^�e������ꤒX�W��"�"�(/�����­w���z����3�Y)�=[����Z7�x�z�>|s�Q�Y��Gv�0��xO:˭e���������^��ү���_����_|8��c�$Y������so(s�����X	���y��`1�&qZ)�~f�[ �[?�C��o��(��<-[?˲�ۡ���1���l�8"ӎb����V.7�"�i�N�\Sa�d��O�S�b���y�rtȝrn�M��z�5S���ud@�ww�
O�S����@�:����/��w����\����E����aX�9��QW���>N��n�]�2X�{�$H�`'1^��cY�7n�e=�m]~�n�l��q�[�ąODʼ���z��g+�k&n��/qCT��=��+ �E58�N-q���:Z��z��)4�I�@[a'8"N�	|+l��=T=��~"���G�F�-|���f��,�Y���*�}7Co7'��[f�N�����nsvv�{�	ey�O�b	_]�`����u����6���#����G�*��?Z�Cp4�L�>��P[ro��͞�����"g�wqb�&�1�g�B���M����e�	���o%2`����A�5���vb�(&���ݎ*t:�2���ު��B�k'S����g�b s���w�GM�@}5,S���/�c�+�k�aֺ*G�]�`�1�-�"N`!>��Aa�u���l�����8�m<�|�ʫy��+3�m1��p7Y�P��5_�n�a����;	�k�8o��K�QqKN�!�H �>}:z��)FH���f/mt�SbO��~�%�$~�q��ϕ�U�\�>`y�V��.����\N�,�R+����'��7���se�x./ /[?�thR�Gʦ�%�;_�v�{�E�И�?���x�?]��A��뗣���Qb�D��f��z�͵�Ç9��)R�i<�1��-WƔ��e�����eX�ɷaͧɸ�o�.���ā�^���辐KV�K�Q�GU]�d=��H@Y�l�a�����<����	��ph���&׶�Vݰ�D��䁚�# D���3��.o+�:s21g8^�Su�+��������G_<ZEқ�h�y��n��.��Ṳk�!` 'KgX����3~�;��rP&��(y���]�(�y��+�^deG��N_�92���d��K<>�ϝO�~xêz����m&m�E�p~q-���0d����y+������}���E&�[]�2�D�+��R�\����S.gX:�� ʷ��	x�D�.���;���VW��"�H�ޭ~���,u�M����g9n8Xw�(a�Ѣ� @��{<�b�5��b�&�t�\�6L"�5�zA�Q�=�ؖlF?>���m+~A�ؙ&�u��l~7��mÞ�	3��y��n�D�@hgU1��&�Z��<��O�۰��o��x��w��v�^g�O�Ȉ�J��7o��u�4����CA�
��occ�k����܃�m�Z�X"a:���V<���o�.�ˆF��aX	T�'�;[WÀ��f��#�s�w/gs��42G5$�&r3`�p�|2�A�ڊ���"W,��rc�F�v�R���S����R� 	�oN;.�HL�сb'�F������>FM�*ڪ8$��D�-;Dc�S�c����D�;��>�%l�.�!vۤ��Q,�yZT��L���8��w*,�m?�Lox���������E5�?�$�[gq���S����^�
�{�|~X��KX)�Z�"B6��It6�	lM���8	�f��'�1<�c:;�gS�>�9�:�f��$�-��b7��� nI���)��H#�-�eN�0$A�Fs�N�S�\��9�\�O⋣�E '���{o�[�!Ĝ�R�����v]��w�0k��l�)���W���D��^�M���Y�FW	��2�ϲ�S��Y�5�߸鯟�ű�r�����/�\��IA����&xwo(�I�wP����o�c���D�E+?�L];�l��|��~� ��H��wܐE<�~�o��GU|:;�y&p��m�vܞ]�VŹ�����B�ƸA���w��B�#�ߛgٚ3˥+���{vӭ��h趰�Hul�u�o�=���(�<L�B����M'R�o2śq�pk���ٮ�.��M�c Nʹ�U�~w)����M��w:��N���?��۸Q�J�y��0���6���#������K��~K�)��s)\��^Ugeu�;��^����|���  �K`�n"�o��!V��5���tTB���f�26;;���7�-��$j��˵���Ԍ���._|���q+Xj_�6����кHt��؎h/�t�M ���	kM��#��6]�G���t�j&.5ϝ��"y).9Q�d+��S2��Q&d�M|BcB�_�3jM�IPg�a}��䍸Q�[�i���v` ��;
�ߑy*UF�u#ORo�Zܥ�W�>v��'Y1��yf4s��������/�8޹�H}�9��<�z��>����:�[��I����� ������Z1���ɫe��+�`♧H�\ì������[�٥�ȗ�9ْ�E���V]=��fh`\���V��i�>Q9�@��m���T���$���    IDAT�"����ݕ/�ԲjyvFj�����3�n���t�[�D����%6?ce��Cq��*A�&βl�0�O�ee}2ܸ:�3ν�#R��L�x:w�\�H[�np�ihMjo�{��7q�����0�b���$UoVІ����a�K�>��۴�o����P߆�N�o��S� B@��<{��=��{��oZ{���q%�2�r��3�l'����u�'W��X'�Y7�u��t��p�-�'��L�w��v�$�����2?���B�pÎ�p�5	.�aF�2��pgQG1��^�|�/�U�f�(3PP��QF�%�������W�%2�2'���O��������7q�8�ծUO"M�{��)sأG��s[)+�pW�[D�X	�C �gw��&Adߵ�TM�6-ADi��v/�-�܍���v��S��)$��DU�79��H�WC��Nc�j�U$��q�G���(/�MK��H�[��55���!
UTO�Dr���h��1�w��ζC�~7;����8v{r�ۣ�U� �э���1ɚQ�_�"t�*a6�%Y�,�r����V}��$ئ_��|�Gɜ��ܪ��ѷ�M�u4���o�^\��(�C�	���/�D-a+s'w � �o�M��?	�8����Ir����␳j��n�r��+���k�D�ܵ���G��C:9v��1ALJ�Sw���QY�C����ݠ��YO�p0~�)��=�&�7;�u�~�����L+����s3�� ��vb�D��&N;��\��E4���
�if�Ik���wʾ�\kgX�1��w>����mJ����V�Z�Y)v:*G~&?��{��ƀ�~������_�P�������d�<��y��	�b�E�Kb�m�D��x��ƿ���U>�W��p��� !"_���6/Ü���e�,W���Q}�#�>��f��s���zsø��DE���E)�H���@fT����xUd�|L˓�Z��W-G¢^�����|��+ض�d|�ʡ�ġs��\���� A{є����p���&%�!�#����E�Ο,7:����i���1�D�w:q��̷�X��K'M�kGcӰf�>�~��C6���kH�v�H`��ʲw9|˥tV2��W����4�_��6,���@棿�+7��~����y���>=����U�7/���?��D�dS���qm��[��p	X�K:��+�'�y8��m��g;��v���!�ng;v��1���,+�Q�R�ɽ%p�77�E���r��Wr��?���f����[<6?tڴ��Y^�C������u��~7��ͷ\[KԊ��,�!��h%�f���=���S��(�W�M��%2�<��F�Vfˊ4ߙ�~"/��_��~"!�d�v���Mf�٣}�]5�ҙ^"�N$��[���o��+�FԈ�h��m�ۘp�屢���+��}&�RUM�,����������`h�rl-?�_������s�K��~��X/��-A�]�-�[��ϕW���Nr���Op ��\[!W7�OmCe���#-��?�����j���n�f���uζK�rleo��S�sc�Z5{�]�Y���*��j�d�Y��w�V8e��n�nW1��(���)����Ĭ��-W��4^e�#�V�{�ز�鎥�NW�u�[�,����=q6�)zYO�ȩ^	pv�3OãL���.�f�Y��w�hr�L��������,/�3o9��6���ܹs���[1J-1�t2��1^���M���N�e5����n�5ͽ�-O�[)�]m>�0�Z�Ú���;T���g7�b���.���_*/��*�a�,CC�/w4^;\�T��𽡂�6$A[7+-&�"�2�� �����K����v���3n�nۃg>��gم�7�8����K��#`Clkh����.�Or��&�؟�;�!$8��;�1����r~��s�l�8u9������K88��
�-�ԌE$�F���s�\<`��U\,aBL�`My���E���b8�\��hÃF�7u��c���\�D'N��� �}�U��]�p�a�v�-���(ko9F�=��R9�om����x�!���X�c�1x6v�{r����N{7)o 3��^�������1�|�g�~�ֺ��{	�I�,'�^s;g�p�U�7׻p�}[	Z&�5О��T���r��8x�����aE�N��X�r�2�k������I����	�㷆:�����L˰<{�K/��<1�ɵU	Z4�����M����	RYo��\[�S��H��>�qƣܻ\v�fź�f�ߺ���ٮm����B��m]2��|"���6��e[|r4���G�˷��0�-G����ə։�pS���6��䕗^�ޗaL�N�~ۮp��|u��0}�c[��ߝ��_�8z淿~���Xݶ���r�6�=�3ܓ~����B���D���_��awۼS�(&d'�2�B��ߍh�m\�v��#�Ry�2_����/��/���8	`��=�Wm��3��2p{;�� �E��;ʈ땜��z��w
�a�躇�X���?7{�k�	gi=K}lK����lN��u֥�}g�JX�q���|��R��[<���N$,�>5�e:1t/h=�MR���Q�y[⒬��/E��<�����N�td�"�c�C�GM��v�K��߸�O2ڍk������%n�P��`*�-�{O훸ٟ�α
}K�vEP��u�vk6Ԋ&��2�͸�N.p�F'�/�Ti��s�e���O~�\�u3��L<�X�������d�"����I�|:!���p�SRo,�t���{���#�7=j���){Kt�:�V��N���#��X��K�Pm�Y�z���]�6��0|n��_Hnz��x5����M=����]:�_l��N�W^y�56>#��+w�"��;eG��~3��t@�eܨC4h'e3<}Mo3,���0m�Th�=����2��.8�n�Ľ���Ĩ}59�e8t�w�}q��L���������x	�Ls�w�y�9��〕C̡��|����=� [�Z�fc������AҰ�`�T�D���x+'ֻ3Q/����0��T���\#�?�+���X4o �>����|���}���5�a�>�\�ݖ�a�����������h��Mp�J���q<���B>|�6�w��8�[�<C��#��y��� G��Wn�Gy�|���C*�@���H�ȗ.��B��'YՇ�&������%!�q�/��;��R�b�����A�*-EوB4���7q�goO���S9۞%�;	���o%0 Aq�)����Fuz��q�&���;�gy�^�I˕s��O�4G���H���V�>��߁����|Cq�R"ϕ� (&O��}{z��E08b�]�)�.��o�^�8*�KW���[ԩH��8	�k�$s��^,$�����x98t�Ӟ����f�� �ND��#��ƅ$T�mgKD7q�p�~ �+�߆!��;�+^�Eы%8��3Uf9�����}��0�]�c�7�R;�"���F#����������C�Y7�w�=������f;$b���y�����g���O�	T���n��7O�Y!�}�.C��+	׳��������9i>V>VOi���l`�8���z����v?�@X�Vgի삯r.܊�u�
��96ػK[�8e���&ǌ�,�jb��K�%4��j�Zը��B�X��ߘ���dM��o<S�s�u!8*�-�?	���QB���7\��	d�M�!(�@I�5pD`!l��`v��-�A�V��?d����/`�_F��h�J�:�=��o��Y[\/�7�b��ǅT�}�����O�K��+Ƞ�Ipz��Й�E�#��7�	{��k��u�����;��|d���z�37pB̂a�۶�J��-�l!w�W4�$w�}s��ծNq�V���F9��7��YBO.�\�4�o��N�V��is��pe�D��/��b������K�CTpqb�[\��� �fń�yVV9�b��� ;��zk�y�X����ҍ^����ٓ���4����y��1.gT1�~�J��
qu(̥�g=Ļ��1[\�4ȁ<r���4�^��1���G��V :�suןmx@d�Yj�7��
d0���u�������E�?^�\�È�*���[��[pm�	8x,���dN'�Vyx��}��i�8�#L�����u�����8Qu�v�����豣�(�A�m��Ia������}�t�ݾ���oqu�pͳ���ie������r�Z� ��~l`r��Z�m:�H��F��.{Ɖ:p]"�k:��P>��R�[�C���<������G9t��pc� FVc!����c�M{�@*��w����pu��Ŏu&��!������S�����8|�KNQ_��1D�@$Y�Q.`�Qmp��P�H�p��IJ��-MP٪C���$x�Nݳ��+��|�vh8��ryul�`�(�$pU���)��`�(&���F������ܩs��+��3��5�U�V,�a�67�
��.I��{��r�?�q�E҄aI�$��s���o��߰��Ω6h*��Fw��������7q�'mJ����o%PN7H�Н�ԙn%��K?�t'��o��rM'���=���|��s9~}�Vs��y�h
N=�PRx6�"|b�@��$$w�C�� ��,�I�A����9�n�v"9�?Z�:Z;�Xy����^�#e���>�l,�l.s���?y�s^���yp��yʀ�b���)[{�|v��M�Y�mN
1:�)�r$�ivr..~z���с���۸�ҝ��2���+�g��d9It���,;��Y�ߖ���+�v��y��v8wG�P��B����;�!;6S���q��[rY+i�V�ڻ|Rl�W���@ɸ��f��%P׹UL �2,>��������������rszZL�Tz��\�̑����d�u�n�lCn%����X�Ȓ�VBi2R�\1@d���uTpX�.�CAf������_�=��n"�om�Cd9��8-�1�ж�f�j�!tdQ��8w���!�)u.�O�+��[Q�.
9��Ӳj9L�7�ަ]T~�Un^�,�w�}�ϕ?���X8h�1(87�pw�\�C1�_�[*gV�Z�	�23q'>$8�������ɟ&������x�]��x^o�SIa���p�.����#]P����b����������nŒ�p�����mY��w0�;��Wy��M��D���I����?��?-W�ވM�n��PH�=��3��1���9�D�]����zH�I}Sh����!�3�X$��g���nq��틤�k�q��� �S�l˙�C7�I���ř�Y43�(���V���P'Q�N}ýu��rzURS�P]�b�"2U�F�7�ˑѣ��k����2�/��"`�+����S	�I���I'��H�h7>��W��t��o]�g����߻�(j���$��
b�����/qGk۫�ݷ�Fzjr*��@>� ���D�rm�����٨�w���Ȧ_��0ߙ^��2�� n�x��������@���Ա3�[�0�����ʑ!�jXG�B��d��|j�*�;&���!W������L'��]�нn��v���9Y>��w��xf�8�gl6F{�˹s��x�<~��r��s�����^��W�"WDQ$��A�l]��
��PE!�ho��{���w��a��q���`�~���p����;��eu� ��=�\��~4I�����WGa����
|*�Hx�7\�껉�꒸}gx�i���3�j^W����}sK��)�엸i���.��Oy��ڳ0֪ܔ��lP �C��N�M�/6Қ���
$���i�y�	J���~������D��W�T�a7��=r����Ѳ:��{���P�ü�~��&�P"d$�W�"�z�I���-c�����9��'k��f	i�z".p���>B~�r��q�Q�NZ:��J�y3gyj~BI� � �W�j_��W�Ӈ�:���w�O��x�|��ϕ+���:��n� ���ݶ*;��Kg��m���5B�8�$\�.��۰ģ�����X'��L�f���X�ż�������{��f����nz$�P�S	��m�#A�!�ފ��C\6��8�Hn��q����U�19�,�i�,D��j�1�?��?���W~�����XH���c9�ti�vq��w%wX{�Z7GE��-OA�Ր��B���å'XY��q^��o$�z-7�|���r���rmu����2���7f�x��N	��8¿r�%T���@��;vŬ�Sm[��E�bI&�Z�Q%D*Vc�l=���_�T^���+�����?U>���R�c���f�GV��Q�����m�"���$��$�H��G���o�mx:����.rɠ����t��:�2w?��J����1�{�=�HA���D�C�×C��3���6"9\x��?�������f�~�q�݌�yq�x˵>�|�	��~����o�	s+�y��������s�|(�^���в'�c�d���	�3�4�Ԡ����v���u��%u��u.�����/��bl
�K���433W�0����r�0��%A�z]rdvv���	U���������gQ��L͔���'������5�E�Cr�3j@ےb��ّ "�hu����K���e<���W�/�x��t�Z��X�	�7�
06;�g�7��͹�scas +CW�)�ݙ����p��;�n�Ww@�p��
_�/�t�A����G7�Э��2�ωc/�xx�z5چ1�3��9��|џ��(q����k�ч���6K����(�����G9�Z�D�6�[foqn���4� ���Q�@u������6�*���B�J����䊇�7��� ��u�2���MN+%����rm�R�m�pV�+P=�+ޑ݈p�h����Ux�����ӣ�f�,3�`1�=�^�/�˭����semv�����~M!��N@�4B'׆���*p��l�)�C3�RȰ|�E�l�SP!R�%�@"����Ы�6�@(�Ǡm&��������{�?��EW'�:;�� n��D���M�ׯ�o�>ӷl/?~�DؖhPW&Y���I�:��]	�^L�q�.�Ѵh�qu�O~�g�@�_��B���rQ��
�����8�����`�:9�8�e�9{r�v�u�v�89���v,�$�5�5;�.���)3��<!�Ц0�BcA��m1-HOi���s���@{�� R������-N�rG�m�^(���*t�k�9���enj��$��K]��n�W_<_Μ8[�������/B����֨1�C2�傰Hx�{w\�?>��ѷ⸎>�>���7Y�����9V��.(�����k1�t��a:[�;����{{�_��F�� ���'��1>�qژ���I���.@��~r[�ɩt�W�~W�.���\�NXݩbz�:1ar�U������+��e�~�B�<�2�|��������=�=�`�eD`�l�GG<{л/����M�£���`Yx��V_�N�k���Ӻr9��tX�EMm�Ё1bূ]�T���U\R��!'/�.����L�Go�o�������3�q�do������<#&���C��,�;i�~�t��&a'1f��~g���δ�[:G�A{lR�Q��3������G��8z1�o���M���#l���Tv�+*�99���M��`)k��h�qXAiu%ʬ�iz;��@|K$	 ��[�t	��9|Y?;�������{��ʅ�O��O��|�|����Ӈ���p��5�U�O_A-ȁ�twޯ��vږX>���[�R�S"���P��z�0����j����xD��Z	Z�n!���'�[�c��hUa�dvy$1slX��D�_�*7�~���w��$6�k}hHʟ���J����[�>f�fѐ�}��}��L+>�	�8�Ig���^�y�����/=v�"�i3ú�    IDAT �U���k�sit�f��E�Nό�7��7q��9*����=0\Ua�"�z�⎎5&[]E 8�����8�k�$��0�m�,���@�5� �@����ջȗ|�5�C ����st8��|=n-'�����_�u������ϣ޷f1�Ef?:v���2�Z�
X�� ��H�؞�N2��٭���v�7��[R����TL��G�:���/Y��%�A!h��c#�GG2k��1�1	��1��0s��ђP�k��8�Z)�_�\�����l�{�'s
:ê�C�[$��wϰ��	�k�a�'�2M����,�g���t��;:*E)�_��,�tҀ�]�5��v�|L�eV�C�l�ݛ��Mܫ�g�8�v@��ɕ�]��z�Jf�k��oSQ7�J�:+nc��6'�9�����o�3�N�z��(2�#��۫���3�~�)綎��^W��k���I�W��g�?Pƹ~�{$��<�h�=�-����5B�\*�=�,�l`qG=)|{�o F$E�Q�_�.T�Zo��h�f�����ǎP�4v�vR��͌-\}��E��l�;m�V���k�[,V=W���s��P��_��r����Ԃ8֗8��z/�]K탸rgRQK�0�w�~�~	_q�8���7��UmȎ�p��0���*T?���e;�vtpqI�J��[{�}���rWo��qnr��~�#)=�Py�W������:�买U q*j�A�' û6V���1,Uߵ��jK�=q�����{*��u�1q]���8�)�1�Xj\^^�ʼ�Q&�p�|�/��q������Q�X
*��'~ۏ��ZъL��dG:mV�RdmU@�#�ڛ��8w�BB��(���3�5*�o%^\[�5�י@�[t�5881bċ���h�	��j�*�`X6�z���Wb���ѳ�y�>���,M"�@��u��4� �0b4���)�#,�Pߞ�&��*��T�Է�ť��N�藿kN���9_�<2���Li���\���ҁ
	����#��#�8���o��M�1���B�@T�B匮 ~�ӟ�=�w���!����R��p��r�^䅿=4�@��	8�@'����N'��|�r��(��	�ᳳ��� �����G~�Gʷ|�{��M�e?ʦ�1�D���̵�r�vc��$�z�v k���F�h�	@]#��#�m5Xyny\�g[i�Wީ��@�|��Z;�Ҙa"�06>`����ȝ�˗����Z�.���W���>,7�7��>^ڳca��.x�Ս�a�a�2B�p�_x��~r�7L���~���S�y&���8�R[��<E��l�oEH�9��]��1�ƚާ��ea�t�o�~��?]}��^����'!}�W| 	��9����V�r �z�(�Z���I�� �hq�S�J��-_������S�
�r�� �E��c�t���Yn��I}������s�S�Ї>T���/��� r�Tg�f��'Cf_Z熭��r��58�������!�@X�ǗW�P�y��u�Um]�(KH+hX�]���u 'J=�x��υ#���jL�jh#��ln�D�k����Y)���	X����K��Ƶ����kat�˽�aC�]�ZtU�:G�g�8z.#r)
�b�ήq"QJx�'����6f�ڜD�针�	�����myvj;^&碘�^�vS����I�,G}w:ӢAi�1�60v��M���n���Y����3����~�޳O�ɾM !"�"���<ATP?}�y~�� *���""��""jD6�����ٓٷ������NuM&<qC|/3V�s��[�N�:u�)�*��@�f̘a x;�Gf^�L1���p��0��*S�*�@)Bj�_=��}2��5�� �@�>��x��pd�����m�s?��O݃�/߇��aG�V[�S�ftӛ�E����d���0٭k{�mm�*ca�����Z-����ڱ]�M�1��W�`[حl�c��k�������]���Q�&!���m�ZI8P��.ߪur_��yb������I�_Ӈ�;�l�k�`m�?IFB�$��aX��i lh�/B\�g��B�p�>}�b����p/��<Nm�lH��Ƞf�H�c�h�g\c�$#��1�X,H}��g����&�S���(ekY*	�aS =F�o���"�}(�^)Z�8�j5r w��ÿ/ @Q�O�eQBCC-�5��&�A��YS'��l����>[�{�J�|��h_w�.v�fN1�f��i���]�ZvS�dqS;�����۰Z���F2'Ys���%�B��T��nR� "�A��t��#:�X�qc�\^����lB�����w˖��e���n�ZQ/fb$x_��̞�p&��$|2�30�g�&ZA}����
ভi��j�жCi���C��7���jy��,^��V`��<`]q3�3c�,# �i8��H�1�Y����Vk���/ܬ��(�SӵЊ�}�Ī�@E���V*��b@ݹVi��7(iQd��M�J�l�J_����>6���K�c0�9
�����>>qƌ�V._��~��t�[Np?�lft2q}�6�DeЏ��aNGsÎlھQ����."�W���+���=����y\)�s?�q��b�䎢��ӭ\�B&`/��L�F���g�*Q�35՘hOL��q{9)~����� SE�o3G��N��6��B;���#<��q^��C<��e�%~צjM
Ħ޲O�n��p�W��
�	�ia�=�Jz"��WHH���H����:/_��-~�b�: 1���P�,篋�s�#����c�$]�Oh0�6��
fqD�U
?��Nު4�5.Ƹb;�N�C��7��l��J�%H�=x=�Cq��ޙu-k_pW}�J�,?s���s���ݼ�{���R9He��)7�]m��ݞs�q[�U��ތxou��8�-p����e�ڠ&t��d<Q�~w��܅��HB|g��8i	�RK䇮v�s1U��9���[�P~>m�P?�����aY�څv`�=��N�I륞�O�����m�R6��4���%nSIgFz�I�`�`��:�5">Iw���� ��:�#�-��	����:�τ�C���/oEKATj�~��x�buS�N5=�F�D�:�dU!���*E�1B�����Ҩ�w$�o���#�.�	i���i2�X�χ�T������^a���+K���MnӺ�n��M��w�[k�Z�0���1����C�/º9��\1-4���II�T#�+�љ�&Θ,=���ս�q߿�F�ZU9��ؠ�E!�~��a�����Zo
�,���.~��扨��6Q=���.�X��-i.J��w�+�!�V�Yh7��M�=�.�!�ɕ>�х�k#��&�MB"̷���я��V<�ʝs�9�U����kj����%*�-��MPs(y��]��'?��?�|��OZGS�őz44��X/���h��o�Q�Vڈ��\�;;�����ۨ֎�v��P1��� `� [��9�Q�c�c�������#���o�{n�*w�'ϳ4k��]����gO��������uR��?g�\7�Q�2 !'�N��ܚֹ���]��ܺe�$�k�� UN��U[�
�&E��-)H���Tn�CŅ_հ�E���H�6�@�Şb�`�ޒD2h�<`����/~�oB�� �;WvP��cI�@t[�R���������l��t"�T�E��ʟI5"�?^�$K���%K0��97�V��QG�.��r9�8��׭J@yp�a���M1��c{�w��i �h�qa�hL�����#�uc���1�/6�0��â')6�<���'bF ��v���s���7�-�~R��*u�C�R�!�s����s��5:����ջ����߹��G��0��(ȵpI��d1�/�v6P��{
�ޒ�(_N� F"����H�Jڂ����q�6UlcE�1%ڏk�p�2��	�½�m�}�INx'\I��̨SFbQe�$ �j�H��N�ظq�o?�s$:y����=�z��e����/��(b7pP�v6;a�V� ����8M��8�]��ֶ���JZ�B�^T��T ��{6#�Ѷ���ѭᘦ,◑�!�_��?�-^3�#�n���#��CHMuX�@�L\�cRN�5�M��5I��I��2i�������X��1u��ݲc}�K��h
���	@2��KV���`p]8�g���"���KPZ=C�+EЫ����(O�*ՀfЇ�c��o�	�38�!��;�b}� ��ə> ~�@�ܧD{�l35#X��0���_<���;���V��^Jrx�2reQ���k��7�p�[���5����W�7vҡ׬_�h��-���/���"���C��l��Vg�ae�o}K�w��vڐ�ЩPn�Wփ�/}�	!4z��5<~�=����A���"�����������,�_���峸�ܧ��Q3`��@E�>���x/<#m~�p����.|x��)���Oؑ�o�?���������^h���ʇx!��h��Ti��$WbS(�9�|��߫�t��o��X�j-�i[D���Ʉ\��p6��N/����ښج�AS�5��w
G��\�B�^﹈�r�* �Q$�Z#3Fu+$�ť-3=�a��X>"L�#��C�gP���~� 2>��wt��<'���yx��t�H�ѱ�m�m�v�#��Joy�7��mra�@�!��^ yr/��o�B\~����|ݩM%BE����:�3�#=�>]��ۛ���Ӱ���< �I<>�r���z�z�Зs�����	�'�n-�y�<)̛����	$(-����pM:2b���2vc��bNb�R���_�����o��ں�8�=����f���_x%|uϚ5˝peU=�]��U��AE��y_܉�KF��p�6��x�w��>(�k�aT�^�A�U|ރ���u���6��H����,��
K�(�u�x��餁�ڋ�X�J��J��r��C�!ߡ�_O���	mae�1V}����O^!.�Ӷ�T�)�[�DV��t����P<{��'�hC�M�P�>y�Ev��ﾯrW\q��1s����[��Ú��[�mU5:��8��r�UϮ];<���tw�;vn}Mm�2F�R�ֹ�J�E#+ڧ�~�F\��fw�A�ʌk����D����)ЎΥp��ꛡ��*t�n�b7C $\���� �͈V����f��"U��a�B��[�6ќ
�Д_�	1�'_iWxy W�����y�锇ϋl����w>! z	��(��6��ƞ�C��w��� ��@эrkVG�4|L���ǋۀ��ߣ��_(���{ 3��4l`)�z��>@����z҉v�rq��s��3 I�XF�)�,z�V,_:�������`j�TxY��c�#7w����6o<��d���h@��߰~�I���U���f���okb2
��0�;�dxC74���}���ǎo��(1����g?�'��C��	�����j��Y�z#�3��"�~�wLLi�l�X�6ګ���P8��0$������h׏��P~�tBk��=��c(�6�x7|H���9�x�
y�+�x��g�P�@��ޡ����Fe$Yz��s���Ez'���/:�K�^�k
��4 N�晪ں<���_������դ���ƍyC[[{�SҢ�9V]���:}��ҧ��.\�����-]���ߦ��v��14J���M���#�^��>�w���\+o�	�ߐ�k�> �D	��sэy)&<;�8Ȧ�_%����-�Y�ٚB)"5b�m``v!?��(8��N2�?(���" ѰbW
�hv�����wf4"��*߭a�o��?�j�3��&m���feo��� ��� ���K���	��v��$/�� �+�o;�dw�g/27��W<�>���j-3(޺�ĮԌ�r⤉9�<���ܴ}{W�x��r�]�m��9��L�tuA� l*͈c�
�u�;����l+dt�YD��^@�ݠ�����M��ڠ
Kk���yp��SR}�,�w̀�:ȏ"+i�;�� ���K��<C�����A�aU���G:�ҳ8�2U�D�	���n�o��)^����!~�P �U��B�֞v�;�	�r�W	����!� ���g(3}����������n�=���Y�����K��!Qv�7�|_��i��v�{3�?^���&%Aa^2�\p[�ZZ�;v�ٽ�}Is��Q�s�H��l��
������>�h�N�u:[PqӒ�$�X@y=�Uq�dƘ�%�Q�0儂��*�k��`q��D���aZGG��#�H ���g"2���sI����u�Z���H�g�a,`l
3Ċ«{����G����TЕ��E9��It/�ɢu֬Y-�@���S�eq�yi�o�)92�"L;����VL��1՟�_�#	��@���o�'芪��D� �pv�ڴ�|m�(���:�Xw�g�w{/��m�l~�Ε5�Ö��C3;�I�#]�H�x����2���ZV^*7�Qinz9�������M.�w�[6o�?4 8ؾ�3�<��pS�Ls�g�v�-RJGY�F�0�v7��~mr0���(_5�"��X���8j��`<3�*O�#��p�ƥ�hX���*��.p�+y� �H�lt��k@!�cpϏ�!m���(��=/Q�0Xi�<��Ƀ4ѫ��8e������w"u���׿����/����g�,�A	��ߡ/�o�N�P���wW�0(=��>��O��|<fc�B?�:�6�����I��)e���s_�Ǚ�g�5kֹ�|����dmg��i 0}���Y3۶�m}$Z�<���QnY��@-֟��wQ��ڪ���2�jV���\�b
\�(ӹ���k)UMp�z�{ӛ�h���Ԡ"4 �)P$�*�N�s�0��������i�Iƞok�H�8hh� �F)mu6�E/
Б�7�k
���xt,���N:��=��i����W�SWD\���AG��l�|�����g+�myNOz�I>�{��&I�{���3'�W�;���#�8�����i_��,}�~xR�A�&� Tږ2��b$��7;���*7m�;>�~�N�p�:����k�ҹ��/o���V14J�=Xm���Ƽ�ql?�|w�UW�~Mn�ܽ}�K_4}����t���1��@[��R����l�䶭��iT1����ǩ�y{�ho�~$R
FGұ�ꗬ2���;l�p��5��O��&O<�[�z�Q�5�AP+ާ����AB�t�8��À ��Q���:���Ω,��-F�w�а�$�ƥ�hd��} @��=y ����8<#�.�	W� �3EB�)�����y�T�Ѓu�ƹ6�_~���ww��wՕW�����HaG�.������|��2�#mP�bEhDl��U���ȍg����>*�=Q�iO>��jm.��p�u�}����B�F�mG?.^�ؔ��򖷺����j���;����W�=��P�G\ۨYA>/3�����ػM>��}�Z�^��~�7>Y�wQ���e������ܨ����\s�Q�{�ױ�y��w��4�c��g�8��FU# $�0�
-vD��������_����V�����PT��0x�@��i:�8af!:�(�ژ�����7H�,������	K�i�{�+&���?:�}�򯻷����_��Wv�4��^{�뮻ζ�i��jX ;���U?�rئb�P��WU|[C��c�%><��M�tc |:�q/u��S^ ˇ#S�;D��>@����裌��r��c�=���/P��V�[���|�?Z=�<^��w��xACQ�b\��\ݘ�/=�賟&�%�����G9.ױue[k[l�dӔ|��( �w�,�Ot��'����u���曭�?աMXg����;42�Y�CP�!:��E5q�|�t⡍���(
��ŉ<���.    IDAT%.�f�G����%Б� �b|A\���'�&�Xo �)_1��3<�Z�����zL�֬Ycu>���ݯ���hqp�s�,H���fР���o� �߁d[�A�E<��C/�6����L�e�.�����ϭdXM�1�#.�ǋ�D����3����=��#������K/�T���;�:���M����f̘ZЦ��� H@����g�Y�mx���;���y���l\�����5+����?���鞆3**�E�C�bR���}���w���E&	�M��j��y���f��F�q��׫$?4�P5�2��K#:�1��s��cu��z	p	������ACU��iO���r>��~�&O�*��lQD���ܪE�2ҭ1^V�D�X,�ʆR�FF���$�����~?+8:��lF�r�n�H�}*�:��a�%e9�$�<�� ����-\�-ƾp�76�\aWT4k/�m�%��LD{QOlߞ���Sqi/��x������\�][����fs�{���I��<���OD�5"$H�&O�T��K>1P�~��[��X֊����_���g��w�x�#���LM,&h4kD5�Q@�l�HTԨ�xB(��;5E��Qg��ޜ�s�w�w���T�$\{��M�qM�4�\�q?]k�V f�� j���#�'Lh���Z�l6��q�[�l-�>{/4C�O<>�tu�
��>����`ĵ:���L�6�\�M�6������%PM�mJ<�Q}�<� �Clk�|ł,���3%PV�V�
%fF"��hW�E���;��$?���ޡ��*N��{��xCפM]!R�3V����np��w�6�5�0H�������96�͛z�ڵ+���/˩׍�I��7i���p�5kW�|��m[#P_�Fcuε,}n@�i ��:���c�ns�Q�.�H,���J�ƯQ����6N$CEC1��kz�, ��x{G��� �iej����R���!��)�t�kש���S��� �Z�\��2`��z�Ϊ5f&" �C�K.�� �*��cI�Ԉ�59�(,�j�~®�&�ŀ�|�Ȱ�2��r�f�@)yT�F	��D���
�;@*vN�!��A͕$�`��q��<a��C�@�tY$C�#��6����GlL�XCm֌K\T[�',W�C��3r�F�-&L���k ��|O�s---���Ǘn؍��cO8���r�-�t(���sPǤ��8��JkQ'������� �dƵt�)��yh7Q�1Ѡ�5k�{�ey�,�'Z��qXV�#�b
%�D:Kj��%�R�S�]���̵�~a�:��r��J���+��j���n��vsO=�4��u˟]a�b���SO��ɛr�'�ʠ�J���nӛ��P07��lJss�V� ���
�ZIn �� p��ʀ���{�����a п��A/W,ā-�}ڇVD�mV.7D%���&�.�\���u�N���ļ�(`O�P(�т=c�@�ȗ��]�:���׃�����'�t��h��x:z��GVJ�U#���8�U���o:��LWϵ�._��~Z��8�"0m4m���\:�Dj�:ₕ3���l�dĚ&Ŷ0ʹ���$���h8:
j�t �y\���n�k=`�uWf�h�C\)�ػ(��1u��P���E����$�$�㘖0�=2T��Fٵ�I��5p�� 5�A@]&��`�g��α�خ��j{����[�� k � ��R��g����͂�z���\J�.����Y�ԋ��} +�I޴ruf�4����f��n�?����c�-�F\ڂ6�p�M�HV�vƫj�(��)t^K9D <I�����b-^��I�
.��y�-Ʊ�2%"DW�$ �`�k��!��Ih�چZ5.�����Phס�]�N$$HS�?jx:DJ[� 
�#�M��E�i�0�����Y�� �5���=�z�f���%��QD���1t�����D`�v0��pHhc��N�(-j�Y�1Px��X��Y7u�4��_�r�/���0��Ǝ������'?$K�I�݊O }�J~�5�-��5����@�FLh�l��%T��}Zp��}�8e�;��jfEzB��5��wҧM
��7�[j�0n�
{��~��6�_��K�ɿ�׶
돯Y��
]%	Ih�����y�鿘�J^�e���p��]j�Ff;������-��M�Ċ�)M�I��]�Ѣ�]6��Fי3�A�ӭ6�.��$^b�t��Ӡ�^	�`���(W���s�6�$�|�E(ZlZR���t ¢�GBj;�:
'�E���O��۸р#`B��� ���>q�JLG!�G�.5�p�#�p9Q^[�T�5Do��c�2XX? 0@�����= N�JE��0����g��ͱn�]���� ��/�-b�4mH{�1��o�f��d�(��k3"$^[l(y23M�>]�GcV��`�x�DM��K����.BQZ�\�(�\`�Fe���W.lٲ�$�R�������U3�l�u]}cT.jeRTZ�Z��h|,3�F��(T������RZ(�t��`�|&L��R���~���M���0=�e�K' ��h %+13�@u7]nu >N�i �CN?�t���-}(8~����<�V$��g���"��Pb_W��C�7�����كrM<�H��1 "6�o��)/�@�'�$ġ����� ���m���6Ȉ��A��[�Eۥ�W3'�����:��9N�1�͊��C���ؠR��I�5U�d,O��w<3n���כ�E^rׯ_���/)BY%��?�����mk�����\���k�xݢlw�ɢ��Ӷ�nk��a�ZnLݦ#.P�ǃ���c-T������f6Ow۶n����H�; ~Ş:m@i�((� ���\s�,�`��MA�+I3�Du�J �)Q�7J�g/�"�N�P���QZ �a_��݄qM���4��*�7ʁO�dJR�'�ڀ�A��ZL�2Q�4KH
���n����OSovq I�R_��.�jm�igX!�)j�3��0��8$���?���)������(�~�d�^���꡶�k�'�� �L̫�]/�R��J�T�֦�\B'B�$��=.���P��+�z�K�m�a̸�wvl+��O��{dk����������G�����/U���Lx��5���>h�W�K�To�^%��Ɓlv�<�j�.�%a�ĩP-�Z{ń:�[G�3�|���[Sʗ�s���/��\�Z�����h���AuZ..W�%]'d����fT�xA6g�~�m@�Դ
�:ƪ���_x��c�ug�u���<��%�?�$��{���c���QQ9ׁ�񌝼s�=�(ã�:�x}�>��Ύ�ݨ�҈׮]�.=�B��H�H�2�~JN�I�����%�a�A�U�1��)�CY3�|����O�W댬6��4 -�V�*����KZӈC�����O�j�:Y�¯�b�T�Wi]���:�oK�}<�7�5�*�>>ߨ��m��=���6+�+���r���m'�,�硕�χ�C�L;h�\�O�+���@�&��9V����+n��K�I�7Zn��`���c�ĢX�L)��EK���.����Tj��9�>����\����D�8քGb��3�ȵ��VJhƃB}YC]�ĐMn�n�ݶ�[���𗀊 8���y�Fu�>ޣx�4<.W�z�ᇭ<�8s�̱��,����B~�E��A�ZҜ�҂]+Td���f$�-7k��K�s���<:�����{�ԋ���Tߓh}��y�0�K�j���r�C�B�p#wYn�>QP�JKg��t�l\9V+�A~1R����v$uPO_n�]��A�#MK�������ܟJ[�=��)�
��w�t�#��Y`a�klH�/��/!/����&���*^{�wݛ��&��J��U0�2l ����;�t�ˇK�X ��qPK�  �C�����Pe�b@��98�%-���w<Pn�!Ϯ�7s�L���'#
e��9�`]����wG[:wĦ��Y,Ԓ%:hs� >��I�Q�yqsjr�y衍A��ǻ@���!�r�O s�����r���sҢ�ob݌-����X�G^�*,� h
�?|� 
�x�� 4���$M8(nN��=t)`# -�yo�	%��yy%~�|)�>�校�(Q(aӦ-�����'� �tI����*)Me��e@��������6Z��i?+Qf$�NKڗ)$"��w�+.���۟��%-ٖ���x;�m�s��Qn���/>!�%�}ƿt:�2c@�=�U7^W<8��AS=@%.�?,(	��|� ���Y�_�$] Gz��u&�!�ǳ���fj�s��@�.3T���hv@2q�%���@�I��!�!Mޡ���J���^�k�i��6R�F!��64��+
6 �u�@��o:�3@`�=PE�lPN(;ׄ�|���i���
p�C������ȼ�=*�lİ���,bаI��t�g�P$�:3^"RN!�Ʒ���N���/I#+"���X^P� hX$@Pz��H�C�uHC������"V���g��E^��ͥ�3��f�pq
� 0A��߀�Ai��F�u�*�;���b�� =q()�!�]���� ��&�O�
� ~�(6~���9Zw�"��-x�C����^��8����klG��B9;ޡ.��@�2V��^Ң����;#�Ϩw,�#q`�Q`QUTI� ⷝգM`3�>�N���`����߻Uk�s+�[54` -T�h�u�Mۼ	@n�YX�[�~;*����\!'~^�4X�p<��g�5!,P�@+�u������}�r�!n�=�k �8`�ts]+�p��Q%���pV�6i�^�-X��~�h_t@[ݩĎ����1*������`�s{�၏n۩(��FY+�o(���u���(p7�t�Xw̴P���Dx�B��� eo�%&]@�~�9���f�(��HCڥ��L���,ΦM�LJ��%�}X �֬^m�ed`Rn�3� �*�;�Ϟ�d��P�4����iaT��gkOt�����m�1$� &	�u��Z����2")�W�Φ�C�k!��֦�	�tmã=��
Y9���Gn,����{�<w���{�9;��qh+F�ZB��cD�v��}�_@��NgD���~kQֹ���H	y�d��j����;���[�l�kٸ� �gH�P�B�	G���ni���a \��k���$�KV��i��>�ܭ�-[�g�>*����%��$PK(��ν z
�̢�{H0��h����=��Z75���1��@(��G?�Qw�܅a�x�7Ņ�By1��;�-*��72;�Y��ʿ���u�]v�{X�6꿇�v�ʐ�2</���}֝w�y�e㝔t�}�)�g����neb��AO\��&��䟐q��wΰ��W��^'�C좶�D�@� > ���������Pn��vQd,�;�F�ަ�[���S����n��V-l[��>�Ԩ���M�ɂ�O2�3(�V���� ��<��Z8_җ:��w�˽��T$��,�Gy�X�F�N�6��m�̰!��O@�O �(�z��S�l*���_�~��IF�Hν�-/��Z�����X����"+�&��� �@Q�Q������Z���}��ƣ�����������S+�'d�7�|����0^�c� WI�Vj��e�Q�a#����tg�}��C<��O>���'-(qBJV�r2U��A��y��J !���X��Td)<E˺3�¨���Z}+JB�����c�] � ��7��K��Ve���;~�K�z�7����b���� �w���<*]f�@D4����5�c3Ė`�N>�++�ɀ���+\ˆ�n�[�w������T�N>���Ԅ{��%Y��gZ�SPo$.Vv�D���AU8�W��Zf���~��!�Q�Nb/�� �`TjK��'��ԓ �o�ov.�7(��-���7��	��	X���7c��in��*v*PR����S�-X�������T��z��bl�u\���3��ܺi�啒,��.W������vȓ�*�f�D��U�F$��Rht���Xr�ع5�N#���2�
���
� �5$>fVӧO����O�4��h��g�c�]G]���OD��%�#M('�� ��a0 Ρ.���0{�"��Sة<���߈zϘ1��J� 4���4y5]>�'��*���5����	�QG���{-HΈG55ː��+`z&�3`$ 5X$$ ��1�eцd���V����~B���S�.8�A'�4	l��f@��d��>��u�ʚ�ubs�u�6�c�9h��e0���E$�~Hh`oX� ?��=���Qg~�ڇ"�(:������i����r^��m8bDՏpaԁ�>�6�[�i�����t: T�5Ā6  ���o>�\9�����($�2*w���b��b�
wđ��H*��(�=���6��#�x�M��}���~��9�����_k[��v��@o ,���x���Pf��~
;���u�;��J�(���'�RuM}�������ʡ�?���x��m� l�`ј���1�@(�"���$`���|c'���*�'��B����jݺ{�<ȏ��/� ���s�.鍗�W�0?'�Ri]r�����	�,��gH[ZZ�y}�k
�>�t)y����y����/KUM��m��,�)���/�(`�Σ�rwvV�(�RbCl�� �e( ��%�;�),
��/��t�����X��J\��Ip�;���C�q�'V��=�N���/����(�9�Am�sf�u�������#�W"��_�t�׸f�(˖=���t�^R���aK&�V��Ϣ�:�3���6�uyf��5
���E�=v��˥74s� XP9~�0�
`��A�s3��L@��eҤj;7���i �@����s��c�I��֜��!�m}��GO�.%i�P/}�Q�#L�1l]{{���?~�>������a��Y�e ��S&ҁ-!P&� [FK+�	�X1q3�L�.�Q6yaDV�/u�6X��f����=z�N4�f �N4����Pp�s_.(��2 ���eQ���ü�։bZ�:h���3r�\%]���z�׼�xnxr �T~Pc|Pm��,qJ��:�Y�ʋ�"���&�-�T6xd��A'cK� Y���C��_�.���喊8��/�mR��SH?�t�Z\D��V�]�ϨdK�2M�ɲe)&����� jz�h�� 0P��ҷ���ϻ׽n�4��
hC�wP\dɲc�)؀{��'Lvλ�G�򁠴��K�kP0S �A:�T�=J�����Yљg���~�;�)'�b��%]�9(�^��w�*y�7����c��)�H����cN��w����-�@-`se2L�PPm��xx�š�o~�ݱr������&��n�M��0 )���CZhb�3F^� dM����W�#`'z��m��D{08�9�S��4i"�����/���c@���H��9����s:VDe����RJ3�����2V�]�ψ��K�MK��,&[�7@`�
���4x]��a? $ �j����S!��}�C2 h��y~`�S�'�m�3 ��<�YCy�� $�	�}�zSV*����a]/y�>	�G:@��;Pmf ����6sDc5X9�0��:�Npo�8 �U�j	��8�{6�Q��\�o��I2e!S�u�go_�͚���r�B��u�P <��q)���R�*H�����v���%����Lx�U�ͻ��|x7H�"�6�b/��_�FMM�ޑ>yF���w�.C����NU���l�ǔ��~ݳ'HM�h%���۫�����r�Hz�G���]?�Np���x����Aq�� �3(0ψ僢c��Vrf�ƍ7���GR�1�L�8��v�H    IDAT7&����2�y?܃�����M����rK�5�<8r�@|�!>� �0;q����r9�}J�z�2BGL�#�:uE"�f�yM���G���I@����6 ��68#�����s|�q���k�I=��qFώa�<�b�]꨸H�(���f��A�M��a-���,�`�`C�Kc� �8��8���e�.��������+g�x�n��[�'+w_^o���W�eg�W�Gz�����d�b1��
-�1 �J��D���()��f�
E�
��{(*T��p> ��/����_l�S�õ�܌��5���\4���т�5z!Pk�4R�((�ɡ��r'L���}��
#�:�����S��V=gqƌmP���ޑ&3��|����v"�Ê
�C�������R.7�dݣܲJ,˩���� ��e��6`� �z�g�����u����v�m�P_n�N��a֬Yn��*��N�6�އ�ت�K0��+�ѧ��W�����s���������t!�� ���Q,�?�Ye�����#�}��,ű��@}�:��� �M07åڈ	����/��L����{�]Jz0
� %�(.0A=s�����~�=����C�����9�'.�q�i��3|���gq�mc|�
s��g�T�0�
�xoX��UU㪙CM[M����}{����;קܜ2�bi��s*U���ŧ�d����R�	��i�1r��F%�[[ӹ�s"��4�8�� `�f���Y�@�=��.;}ޱ�b,
j��i������m� �
o�Q����o~�'Mo�aM���U�V�ռ�sd��*^�ޥ��L�ރ�6m�`,�\!�V��B���ꡛ���r�3��h&��{� ���Jp�K��qݸK(AY����d|�AE���H������v~����ͻ8MFz��I"h�Э^��s�a;�l�N �,6?���L�ì �vX|:�ޤ�D9ɏ2�`�r��x�y@M��C�>�F��O��Jԯ�%R�K92Z*5F����r�?��Rp7'$��PƅS5�  P@��*I?X����:=���E��ɍ�r��!��/��s�央���������Zy[z�j��轐'�JLF�-�>��������7q����ex��V-�\�6r�f@ןH!& r)��M���F)�kd�U,��IPP��/����a�sB0�7��?���N�c�9w��S�����:m��#���~^Rxf��'P߆����|�m��T�����A~�,|'�� )UyP{@��4Zo�p~D�lJq%�)��6�T$Y����m���.F�H��{��M�:g����7j����+iȾRȨ(S	 ���&��5�^owK]�v�}w;�]���i�C��y���FM:% �3j�E�
�<H<�J��$����}>�v	�kn�s(���9���=�k嵯�&�m�( M\Ր%ff�x�H<�L��u�bq[���I��W?�w�
�E��J��H<p��;(�Oj�}>��zx�׭[�+y6σL��X` ��	��7���N'ع�0i�'����^�V_� j�q?�P����q�v�[[��Ӊb��,rB��u��%֡"�L�~���6ʆ�I`ة$����x��'��?�+��`7ؒ�?�e;>�+��b����WG�J06P�z� AG�A�uO���Y�Qhv&���;�p�u�>�Ry_�e�&�enN)�Ydq�4@"^����G#����%����n;(=~�V H�X��
~���.���,��?�pw�G�3G���@X���}�{F�;��tD��')iB]aCB� ���oE��}���n��`�1�� z�D�U�7-���B\���s�Fp�_�$��E��~�'�C ��W|���zM�<���o�E���/��G����*9��=�AP�[����tn�5�Ɗ��F�mSm�i��-J��h	b1�9������Sx�.�f�x6U(i�ғ< ��N�1ʾc�}�<ŚT�pCg��0J�Mח�=��A0 x0���;��,��PrO����p-�Z$*nWW���y�<Ɔh���Ve�8�4��X
xl���q�Ȳ� "��T;���zXy���ܿ��H½�W�34�dJ�Hm!y�8�=�o���Q	�f�+E��82T��j��"
��=؁�@ƂL���5Y��g���K+vZ�� v�O����=�K�`����t���Eb<Qc:)X���X�{ޝM�I0�'"�D�W� �HL������Z�+Gj�_A��'©�F��#�gsz��� �`[B���=)br���b�|��^�nk�]�O�X�}u䳎���P�^�"H%��P�`^���l����@�Ȱ9��=�y���?���o���x�)>a����w�ml�� �� b&``J�)��.�=��{�w@�E��h�fMW�YY�4�t��	���C�<n|���!�KN@�(� ��7΂�="¨��S�dl�1!bE�5����٧"������ )"�^D|�z�:�æK��6�Z�;񤷺3���|N�n�4�d���o~�D�u0*���|b:�<�ʒ�)��+j����J�`	� 1�������à�:�rhu�7��B���0��ފ)�Q��_��Q�!��"�����������P3> �Xr� u|��_�>���X���E���_��TR�/_�V˘ �$�{��d%���x?Ҥ� �|��� ڂ������|���皼�;!@�0�`��w����vC���{SC8�ܥ�2�¨�@!33W���C3� 0P^
�*�>5 �x��ܹ.)����o��g�=c:�����g���ȇݏ~|��#uڪ?P��˔DR���PZ4�2b/����-�m�`z�a�߸�t�!*;�2]�B����}��K�}��p_>����+w1x 8u" l��:��1�KxR�)�}��C~�U�/UG�=���� ���xh�y��^�O"A�"/��� ���k�UW]���PMT[���<p�ZFܬY�L.���,^����	u�U�;q�̙c�O��)����ɓ����a�\F�N^,|��./�(X���{���~� .��R����b21aTR�͛'絃#��-Q����Ȝa�+np �E$�ڜE)��2��x\��)İ=:� �� �/��U��I��@ ��cG��QXʄ/p�_M^�Cz�U���=�'��)7i�<���\PtS�1��|�,��#(�JpK�[�+���K4� � 
((�� ��@�~�[�j`�3{�[��<;�:PȦqM:�}��6`�o&�ːg 6y�>��;z�\y�<-l��j�b�\�QV�y���_kG?i	�����=$@�E��wKd�3ْ�47�y|�ˀ�e -W@��X �"9�+T�@@	P8e���W���u������Z��w�o�p�Q턬o��#�6?)X� #��a 1{�7���<�<#j ���ǥ�W�
F�L�B��d4���%�F�>�T�V�6}�s��@���G#�#]Cq�I	v��� "�w4��2�����׿6�>�ܪ�N_������7$1��h6i�dY�<����y�C���E�Т8�o,yB���A���P77�4�5Y_^�u��R��V�j��0X(�^r��3�$F�#崄&m0R#'�Bpۙ���NG@9��w��QP���b\���\Š�nYڰ#�+m?΢D{�Z֭qW\q�m� ��%Y\'�~�NF����h@�� -�bO)��	f��k�� ��9���(�ǈx���l��MF�I�4JJ�r30@U��@�5�C�7�U��s���ߡ�sT2~
	w��(�RM����L�4��f�mSE @M0Ê �`�P��8�?����7�k|�X �����J ���%�m $o�-G(9��������{�x�bs��q�y��,���~�ӟ�Ye�]�~J,3ԝ5 y��Wyi�J�U��
�#:Hؐ�J�e���_G����Sj�����&H��\A�?� ��ȗqd��!�e��@�
?�;T����F͗�� �8q�Qq�p����G�1!c�$b<��y�)wU�9�dNI���7h��j7t�[��1�-�}{�vw����.���::P�4X��؏��zP9�W�A�_����x*�M��۴|^)�Īd��吐�aR�^��BJ�������}9���\9�e� 0��Q9��v��x�8�u�򖷘��I'��6h�/��3��#Pl�Ǖĕ���	Py����;�^z������w���E���Or�i刉�&M0��>8��#7�%6��а+�	&��E3p��7�{D ���EF]hv�ڏ�09��K�s$~X�q?���<<n��`SPl���(J?V�6Y-,�daw��xPu�3hx�4����M�[B|���̮_ߢA�^JW�R��"����o���9��Ӄ�׃��d��z���H����ϖ"^ڮ4�X���0*)���zmF�n�'P��n v"�y�t���dܘF����N�����Κ5��	�2(ؕ������%�Okq�H㩧�rϯi�"u��ڨ��.�E^�<��r�)�u�}��ݯp���o��Zm��R��+/� '��R�4pٝ�+��r]]>&Ǵ#&�Jpo�V�O�Q�K$������\Tږ�ڂemW���=x�*�'ݑ�ι����^�׆/�M��dQ�}L�@Vi j����Vz���㮷+�>t���S�~�uw��"�3�p�v�����m0��e�0�`]�'�v���)�LJ�Ȭ��J0Lf��o*�ŒD�N��L�$)ݪ��8�]Y�d�;۶��0���ޠ(UL�~��9�sg�)½��p�2˨�Ă�%���;+`��B��x���ũ�K��&����������"�=������xu%-L��ȏ`���Ǐo���	�M|t��|� ����@�=��<�m�l���D��g�zxgW��:pO���FS/r�L�\('d���et:�ۀ * A�l�e=,�@��K��K��J��q�������e�N##����7�!��k\���ɛ���뤴-[����֚4�<���Nw�]w�^#�9����{��$#c��z��d��l��tv�[�h3Z}�~zqG��]�-�-K�5RNE��VI�c$�u��j��t�$�G�O����nE�fW��Nω�'ϡ���PIuȦs:����KX��caZQ����[����T�k_����"TT�LZ��s�����]w�Ҩ9���
l��j1�f���t%���:[�º���ڀY	�f*���/�"ۚ�4�s������ۋ���Q�͛�����������w^d� Q��. ����η�==�A*�A0)|����NV\rl�?0��@��ء��ץj���Z9�!-Ψ���eu�:x���f�2��4F�6	����D����?��ΙG�����@�Im�)b�$�����c~�F���D��=<��>���_�!Kl�$ئ�Uq���!�30��p�d yH�g|X�A�y���{��ܩ�u��`(����	�	��
�>����<�#��Y޴�o"�M�6����m�c���G|h�6�[Le�]��#�x�nxpcY�P^�[rv-j��6�["I� Y~K�""�ۨ�vu͉L��>��}�1ڃR��Ϝƫǡݺ#��搠Lw���5�����;44��^���y9���{��,��ig2#�Tݫ�j��(� ������wާM��6��?�cF��]9���MD���0�LŢU#���$Sq��)=�*��g�J�#GDƐTTŉ�b��v�MV�K��(g�>۝��[�]�����.[�����i�2�S`{����C�PZtLP�x���M(e�v+�;�=���7i�4��B�o��;��xagV^{ݺu�!��a�抂�1N�	�(�d�	�����E?��6w�7ۂ�����9e#UB��oA[�|]*�j�N���xD6Ŧ���N<1a��[��u��~�S*�� `����d�P���^�	���<+��E�<���lP��:�v�W�8���;��Gf+��W�O\��u�Yn��yn����c�u��DVi��U�쫁ǢW�M�x�I"|8�P�/�%1�C�Ć����L��zW��fiE��m�\i��|�N
���(w��<E��Ɂ*0�7����$��_��W����A�9��j��vj7�{�ᇛ�5���܁j���<x؆g�%��'�x����Ysܷ��-W%������� �o��-���ƫ��=[�9�����,1Pq��D��P}ṙ��8o�������u�܈�RG���e%�<a�ڶ�� ��v05�3�s`>����k��.�:��G��jɣ���'�x�]{�5bn5pV���.�HMM���Y N���I�y��2��<��3,�s˴-��C��"6�*�|-n�<Xi���8��*�f�2@p���1�侴K�i�%C�t@N_��F�#(�R�-y�h��W �ȕ ���9�4��z$� <+���v4��O��S�)'�͜���u����`��G�Zs�5� ����<��'+��bTP"�a��ꫯv|�!�5ig����@e�kN
V���J��d%�ā'Ѫ"j�?�!pbH�Sn�x�3b[�v4J���^G+��+)Z��I}D�<����N-����4�ۛ��f��Y\�yƙ����=��f���}��Da�lX
���HW��J��Gu�Q^�5�9�2���v���)�O�	��W��v��6v��d�<�/��^�,�a�FL����hR��u N4�Hź�������V��W%%Q�,����kT�6 �Tn�2�Y8r~#@`��z�9�8�(�;�\���w�{F�0u�]c�V�7�1�q����x�������w�_~����Ns�Y⹱��w�}L�kì�A�ƍkl	�ܤ��C :��UZ߅cK��3D�1��r��n�=/?�����QJ���'WN�X�BE��y���C���hz�+;��$��5����-�P�u�ofc˜3�<˵i�v�Drx��EÕW~��a����Xޠ�A�Ix�e��o��s�=��ħN���XHH���{6�J��dU���p�qΖ��ճ[�bMT�WR��f��^�u�Bk���.l�?*���ԇ��_�JW�uؠcz�:C�q��w��3�">��;�x3F8��%^�Y�R�&H3n��FY7�"��gFJ���/h \�^��W�Q	��Γ�p�6c ���R���g?��QO�)3;�������L�H4VҰ��P�}�`C��ŋG�٣��'�ږf�̍ʻd��L��Udق���E@F/C=��%�@�˲�߼������|���w ��&
�����E�v�Ĺ�R��㠫MhsG�'�X�5ԍuw�u���W�po��7��u���Z�x�gW>o3I��(�m7�%�ں��xB�`�s��|��L���z�r���_�E�#5�4���-#�x2'&�ɘt�����a��w�n{��A�*����΁B� ��� '.l���z�灳}.�Bг1�]��l�d�yg{�(��� �/���'L�5O�΀op7�p���n�r̙;�]t�E��s�������u�v�$۲f�x�:�ր^��(#�0ȏ@���2����l�U�Tã���������Bp�ism6VG#%����~��%�\:<#�a���W�� V� ����>QO�shp0H�o٪���J���?c�N;�Ĕ���Ci�0����f\�����=���n�����`N6�o�$&}n}�����g\�FR��2��'aP�'n(๽��zl�ʈxH�ע�T,ǤӞ��)h,�\�Ī:"��Jp�ߝ�����RI6�t<����7T �lap A� |�J�X    IDAT �/}�E'*<�j��=)�W(:���\���fhx�4��[��^{.p˞~Z��:���%��K�R��W �.�T�^����?������(0�G�K]mM���V~"�=e'��C��pWWWe�\H�k0ީr$�.E�Z���0*��hM��3#=�m�<�έ:�`S���7�̀�ā�#��ꐤ��z�H�Հ�+^NԳ��^[��A�⮮ќ����	���wP}0-TEȉ�K�ɀι;�h
�� Z@�����m
E��n�f
U�����m�P>��ͯ8N2m�SbK��k��:��}��k�L�+j�s��;*���m�O(����JP��g Sw�uD��,9r��[l}�]W�t2����>W|r�d��i&������Q�-
���#}@K�Ȫ`�Ƣ��SNr���g�#߶�E:.���Rռ��K���X��6Uq Ȥ̼B �ؗ*�Q�蠺c\�)�e#K�W�����,�4�^��
   �^��%�Q]Se�.`d L���}r�v��߶�X�#�C?��9vO�����e��R[�C�D���G^�>��=���s>��&�����%`w�w)mY���� O�:ո��$�e�-Ly[��5�$�_T^�JD�P�H�":f���F|d�Q	�������6)^!���PR� �
`r��*,2m�Љ��Vt{�O����
d?D*�F�Y��@O�֘� j�}[�=K	�d��mh�f���w��5E�{{���~v�]�*�(=R��.��7���}�B��a}!㉼�#����#bxa\G%�{z&�Jݫ�>�{D�j�
*ᯁ���5K	8�?���G�O����x�ݴxh�1t�C�O��7*�����d��b]�.��꼤8�d�_����ϓ�b�5߹�=�j� ��X\�/WJ�-�0*�I�0",��"~�"wm�5�lQ�[�dA��m���(G;Ӊ�u���}�T�o��v(�R�P�p`9�~� *�(|�:E�a{[ �k��n��y�,�p�H�{����j�|挙���	b/Z��&���m؊���\}B�B��p���p�������D	x��x���|��|B�,!�Q=�aB�5�X��∣ޣpA�"=�MD�R�X!&�-E��|�H��NQ�:p	��[�n�֢��f���p|�BXW�~�Zyb�W�d�;O
O3f4�$�o���U^F`dA*��z˛�e��#�&Y����6�p� �f�� ����)/��<5�`--�k��-+�m�����@���h�>emK��bI#�n�b<k��#��\���Wv�0
�]WΥDBc�y���$l�- 0@���?��Sm ��T�������1�EC��矅$O��8�v�-[ni� ��/`��-�k�j**�Gy��K��a�`��=��?,���~�Iw�]w��+N:�t��ծ�u���M���zK�هن4�5�����Ŵ�#ENX@�DҒr$�b���ҕ]ݣ�Kd��G�X|ugGgj	�� ,�l DA�)�HV��
���>c��'���������vy>�� Jb:���(�?	�CI�?雯o�������ڵ����vBZB3˥_��ť��o��M��\x�%��/\�A5Fik!��a`�IT�Z�q�0X����$�B��T90��{�0B���NTNVf���>��PQe� P�+!HF  2n���=V�
h�����i�l�/7MM����x���S�E&�,,�5H�ee�9���PU!�Hl�ڵkm�g@b�U+WH��j�Y���!^��l0�����M�J�����BiC�	<��i��{<�'$��+�r<�!���t��0*�].W����
���`���H ����
O�>7� �W[#����Ǐ�`��p�;��8��)�`Q3V������ g�˳ �h����cB7E����N�'�|ܽ�q�ۦ�(OR�,o`�pȃyT�AI��N �a��@ⷼ^u�;�P^�dI����6��=ɷQD�I�SH=T:�Ѐ� � �~�1`Y����D���^w��6e�[�f�tLnv���&��B���vx��`@v��C8w� ������9*��:���w����̠�XD���y��?ވ��	�)+�����������%�Ή
Ҙ�೬�93����	��r밺��i�bNC���R��xa|{���7c�$���Iz��9�Z\WG����ϚYF	_��W�;O}�9��?�,�$B���\^��;�z�������C�VEnDO��I>>k��֥H�X�-���5JLR�Vq���W)�qQ�I	�A�`����w3�f6"����LjG*��D^*�LJ��u�{ڴ���֧�W�Q(t�;���HI��~��3�k'ˁ�M7�d�ϐK��+_��[�j�m�j�'�S���抁S�8<�c���X�����Ͽ�����c�<�#��VF�LZܣ��7l����!����q�/.��u�Yc������5aԁ;��Z(�38�7F�5⇽~���NlE�:�~��6/j�V �wJ[�Ȥ��Dj�6�� ؂��OMZ�nI�PxB�;��ʎ)]�]��>V'������Z�v�`�}� x���� c� �0H������d�5�M�T���rz�܈�Ĉ�H �K]L[0����1��oѱ��eB��O�^� 8��$ ����d�	���X�[�#�wJ:��GG<�@�B�|�_�e�=���҇gl���I�SO-s��|�r�����WK|�x(JawI��@�\ ^�8~0���&�^��������.��bm�0�G�lD�V��;"P���,��5]��9\tq^,Q54�B����0��zV�<Z_�M��X�3�M&-9�E�/}�2R@>i�d�+��pw�_0�w�j�������;L�5�HR���R�ɓ��N'�9��a��PZ_�hZ�����˟��[����U� = �+�D���*hs>���W3e��R_]}�vF����Ė/_.n�(��v*tDr+n��	���v�g����S�W�F'�Ǝ�wR����y�m)��,������2�3�=��$b59���O/�0<<_u�{z��ģԛ�r��Xr�d2�)[� �$����P�ԒE\WW�{����<q�D㛡� �<�Pf�#�8��}�<� P������X�2��T��n�͞1h(#�D�-�}��J���#Ik��Kdzr�����R>Z[;��;[մ������n�xi�-X�t!� �S����K�5p���/��%��д�iӦUikmm���j���:M��������;���H}~���'F��I��hYs}1��b��Fr��&[j΢�1�.h�!Y(E�3��HT��ڷ%J�h��ݚ�d��մ;�ر}��Ha�<`6�S����렣�u�ف���G:�mj'�@��g �k�q�s�"Ӡ�o �I( �Xe�����^:"8�� .��	����4Pa,�E9�/$ZdJc�|�0��ߋ�x�K���.�ރ-	&�s.����	0/XZ�+�����-ֵ�u,�0cƪ��{L�Z*56��*�&L㸆��]9�ɕF�b,���)�E92k�>:�-�(F��h)Z,um��j!6_��do)2�M工]��N������L��4���6�reK����Q��K��������6�4�Iɪ�"��I�a�H�8�*)X.�uu�|Ok�:^��R�ڀ蕓�Bv SǙ.�BNjrZ�E�E�S�G2����ܪζ���J�\���6։���H����	�C����/O 0 pf(F�� ����I��28|��OVD�H. ,:( 0�R���-Gq��2Q��T}܄q2W�Ii%���Y�:yse���%�	�b�.y00��.�s��M�ԋ:�qݫiH�^�d�ɾ��f�ŞX"9X��z'�tQ���II��"A1���"b�
b��IR��~����b��:]9����<����3��L��*_̯�<����n���C��j�ͷ�?�����/�u���x������T$�O_w�Q�xdL��;�l\?`�%۵V:�¢���v��&W}���޾�v��<�eiF([H൰�&�^��b�!�l?ƻ6`֬��^���
c%,@a�����H�:Ǜ�������5#�[����*�:�ԩS�NUQ<�2���f�8@=tY�G�ճ{6�@2X�fx!�3&K��1 ��wٝ�^9�L,ɨ,Ϙ��y���`Io��r�<��\���j0�i�l%�A�,��d�Rn�����~�G�׽������%=V��l�rC��(e����?x0s�ո���W2����5�!������O��W�n�<�Kc^�W��ԳJ�����ҧ�N���{�{gwe}ue���{�ޓ�޹ra�����k�o��{���ǟ���o{�;~$�~L�����>�03������W�f�F^�v��3�7�����Np0�D�Yx�T�B4��R���	�m�S�N�2�A�uu c�g:S�;�B!�⊩�ػKj/m�݃��	�k�W����a ɿ�7�F6�����S�xO�L\�O׶��]_����.K���ͧ��{�~������o��L��#a��sr���A��{��*����Gԉ���Gg�����EX L�YyF,�����ԭr�����l|�<��U�C��O��4rG|7��Çv33|aucm�����pbym�On���>�zv����?x��Gn��ޓ�W&������<���x+S�^�g~���W>g�Z�gs������qi����s)z7�{�H�Ă�xn6�n�,�c(̍��`!d�"���U�3��/��o��L�
D��`ZK�)&3����~��"!w�E���΍	�$���������ۓF������w��\V=��X]XW�g=�Y�O��O���7}�7��Q�q�1L���!�<]�gTou.���ׯ�i���3�z�6�h1�����i�>����s�v���<G�-�w��jYc�{n]4�����3S�ֶ7ߟ�y��������Cǟ��C�����2���DV��Hq�K�No}Fv�y���Sw�̎��DR/L7�/��D�/&��:�b6�~�U+�a����ǃ��Pq���O�;�R��.�e��N�C��75૿���Lw<'��*���E��QgP��7|�7����������g6�	P�g�:D]�jF��Hy�t�������������u��G�o��p���aR��]���7u#:r��5|���:�bp�ŬE�z������mu��0F�)G\|M�e51�g��m����3���o[�3/�랻���ͷg�^�s=>��=�O����������/���z��>|`!��r����;T� I��w��t)��#&��Or!;H��Lg���dt�٬��q8B�D�`Vя�2IKj#:�C0&�lW�"U�T�N��O[�BMZ��ݭ`g�+}7n�t_�z��{�Sy��]�Ƥ�Ν���7���_[�8R��US�����V�!�j�`"���o��᫾�k
�����L�	��7�����8Ĝ����gŽ�/���d��w;a����dZR��x��eSc����kX>������=��c,��e-�L< �����SK�/�˶O��?~��#7���>�߹}��F:�� �@����0w�7�n�����寞���ԕ�g����9�ըU��K�d��[���b<�q7��}�6E�q�+B�Q]�i��t�ē��(�܉�Ӌ�P%�:��]Ҏ��n��<Iu���OD������|�v[�k�s��w4.��g�X�q_6������B4㊇Y<;Ռ�ˑ#7�����,�J�.���շHkV�ƭ����+����о�M�p��O޹��ңw`R'��r��ā���3^��hc�ӧ��?���x���?�1��dm���ý�ؿ�����{M�bn��N��~ڥ3g��?w!���# �6KZ"*�
�ƶ���9�T�B��;K���A>� �"C@�w^��S���b�j��Dhy�fR��H��oٮ�7$GD���,��Q��vT&:��$�W��e�{ߜu��$Tҧ�t/2J�q��+��j�H���F�ǳ�ál�Y�@}T�������c�>�|1qMjh�)w%�U�:13���w�޳z��X�g#S6��L�*�[�7��� �w��מ��~�OT�Ld��"����h��d3�&��˱)b�Q��r|]R畩;����/�����S���O�m�|��<<�������0|��ӟ~iz���o�\������?�cͨ@G$yf-�q�K�Z��C�|�h�?�ư���/)�FD��|$�W����V��C��nx�w�S*�0��`�%_�(ґ�&W��]�ӧ��x ��ߪ�ģ���W~�`��>��������8����2��˦��F-�����|���k��kU���\0�9��J"+�[�n'�QSTM����u��W�2��O����4�������)=]�[�}��* 
p�^ރwf��OV��fvh�!�ď}qgys�O�f���>r��ҍ|8HO��c&�����|��.�^�ҍ��ϟ�\�5{I�ؿc+��h� ��JAߐY�a6��pQ��Z��$�3d��^$��3�l$'d��J��T�+m{���f:3�i��]HL�Uy����^>�'RK�����NĢ=��|6�l�c+G��XC~$֍/��/�e���%/��bd̪�$���U񅬆��c
| 5����V�=)WL�Fz��ɜ�v2:h, {&�1f�\Iaeß���uBS��ta�\��q�L��oA�ɿޥ�9ݪ��$���v�2Ѻ늩{��U����҇u��/-uI��u��v!+��8p��FއƛQ�&Z��X�,������}��Ɇ��0�ߖ���r��G�6�"�E>���W<e���?�Z9��O�8�"ڎ�{
Ѻsā���QK� ���B :e�뾈�u���� <��ż�!����K����K��Y@���C�I�Kc���7��~����S�F�	$=��bz'���!P�Yx@/�c�����L�R�^����^�����ۅ����۠W���V�^�՞�U�JH���R�s�+ߙ��{x��-��<]��&$���|U��$Iǳ�z�Y�2F*���#�mrh~~vcb~�������ڔ�UE~������b~ߞ��W~����^[�x㩓��`�XWX�T	����V���vk*��׆ i��k��0o���֦�+$�N�����e�\za!oļ�������W�z�^�`
֒^7k%�C�>��R!��7d�8Y_X4�k�8����eԱSgN� �0�`
S�/=7�I��߈��p滼{��꩗LГ���;�*�w~p-��4*��+8���iq����^~%�o�kKs�z^&�X�b�Z?t뭟~�����>z�����w�N�ϋ��|��֗ޱt`�;Ο~��# r �Iӆ0�O5
y�!�*�\�#H,�.�p���+�t�.�K��8�}��l.�Yߣ�\!T�����o�3�]��|]����l��ggx�6�w!���<Lа�aYN�n)��m̷���K7M:�.�TnjU��G�H<�G���ޘ�6^ة��V�����D��+������*�phR�������N���Rz�v[���S�J�P���/�6?{h�����QM�|̘��g<�kN����;!�� j@7�QsU,̑z�@��~D�o��W$J���Wi�����Y���&/i��iDH^tu����C^D�W��ؤ�P��nԈ�&eC���1Q�9�}+u�٪�F�b��=��R�t�+9�4J��w��#7d�Υ��rąem�\T���.:�1&{cd�jvz�'0Ի��`���װG�
�����z�c�!���T&5�Z�v����aΡ���A��[��QgzV��qYp�!/�S�
F9$��_$/g�onj�ݙ�[��6~>ƈQ��œ��1��g�����y蹵}A��Pk���P�{�p��|�
���uDt��Q���
����M�;�i Z�(    IDAT�A���z��Ȇ�$����J|���r��<��~�JJ���w��T����ʵ"G�����5n�6ÉI�:�ݷ���:^֕G�Q�]�����R���|�����/�o���U�����p��{5sv:��a��Io�y���v�1�hf\�^��鹩����55�I�'�$�>&�}��Ϻs��cߟ���ni�R�9��u��{e�G��8.i�M��ّ[�tŝq��i���l+MbW���k��"�����Q��J�Ew���mq\%F4qH��0��6�D|R��b�����+8��//s������e1_``*4Ѕ��8T��Wӝ��$t<�����_%���dV�[ƣk���ge�O�j\���GȢ�<-��~י|���~2UT���V�-d���&p�A\i�+[����ixe?5�rg{cnwfϹac���6e��D�����G�.^~S/�q~�;��f%{�	T�.	 ����p��&qB@i;"E���tfw�w?�;�����g/��?]�5¶�:L�)�Y+�����K��tkR��NiH�Z�������pI���]:eˣױ�������4B7��o���o���=2K��ǵa/��_�>�wX�������Ckߥ'0�(��峇8A�<�t-�>_��>z���{����?�l��E7�U7�RKn�F� �WƳ�{'N}+a�/[%1is�W������S�x^9N<�z���x�ίK�e�.ť�^7N�ҜU��!�t/I��Ҁ�RU�Ґ���t�M3��}��W�u��O���)#ϥς�b��!ӣ|{�������M`(sq��.��ΕOz��oD7������������|T�2UL�|`wSz�C��D��HeB�D����j�=��"�dƲ��#�%W�������/6V_nj]�p�h<K�5D^y'����<��Gs߉wm^��o����w��w�(N'��n����0��4=�o���u���¤������?~�������p~�`l�Wur�)ӕO����^�t��`�^���^�w�o��;�V'sgcF�{��\Z�A]����=C93;w����ot���uC�EܦZt�_AT��`�IZ-4X�v="��b녺e�~ @>���y׃wtY��`!]�|U�k'-�밺�!��i����Ο^��ʾx`xA��_@�_+�ʧ��I�OX����
BX������y9�<��奣��������o~�!q�K���в;����g�l)+���`+��J�ȧD�6s���~ol!n�t���Jp���粠U�������&�o@���7�ẙ;@lB�[ٚ`:�P ���u�"W(/n�<C|W�C>���G._z:��8�*XZYWผ�In��iy��c�������~�
~k
�Tp���T���_O���
�t؞(�eX�m��v��zW̗:=02�:�ۜ������I��No�@>�D+�.Nm�f��I���J}�1^�N\�����a}{����ŻS�Gt�^��j�[��|Tq�_˲�n8��xTP�F����Ō�B]�.V
�#f��t���g�]�B����ECZ�m���&I+�|��fr/���t�K�$��;���D�~$E�)kE���X�Ȋ��F ��2���K�$��a����^a�n�zW)1�7����a*o���O�ޣeyU�'��U�x����l�ٟ���m��2�e[�c'ZG~�3��~�r�ک�d�R[a0���][w
[�5llm!-�OV�e�#u�"�ɐ�s�{�O�$�u��qM�^��	]���Y����[m���3�8rլ#\����R��!@Iki�$�������/smp4�,Ď��oq��v�{�2�n���'ʣ�8�(#�5䤪t�6�+y���z��(���0����c#f�7y����i�{a�\��Bُd����'}�'�5�B$�ox���t�-�Ui�~{(��])[�w
���#���Rv���+��
�v����K��ܸ�a8������2���yt��<�,�+�?ȮB\1�HH�BР�������X�;QZ-���1+n>U�ѻ˙]s#N+3�b��E�� ��	-�����S����*n"y�ǳ��ӞG�I:娑 ������>W\>���c�	���*��Cj7f��
��Ԅ���ٟ7<�YώE&[��-��ٟ�%�4�C��U����?��/�Ҕ35|K\~9����邋N-�_�|HyW��\b���'S�痟��/�;��=����u���{� �<Q��^AxG���W$w#gϧ"��H�C/�?c"i�u���L�zz�����ǻg�����Ov��Fx�l*��\O�g��`e�k�ӌ��^�h��HZ�z�)�;��ӑI�<�7&=�0����o�NX_U4r8,;���re|����Oy�𲗼�xA>�eU!��tT_&o��{�bh�ǭ����w�v��<=w�0\"���$x���ލ������ B���s�v��Y��X�߉Ț&�tˍ�*���@�˱�D-;������t����F����� �'`R3��-Sl-JqE�*�Z�^�	2'R�PD�UR�Ce�Q�'{w1F�[�3�[g"׺/"��K�[A�).���u�[?�{�<�7��I�G��+��`+�_;�/��78��-~�"e[)c�n�")W�B��tɊ(�O>�;}����9ab-�3o�M����l5��j�疲�KV-e3���f�c�����d��ȅ=sSi�ᡝll������le]ힽ{v7&��H�'���q�φ [(�iE�0g&�;1��A����K6Y>ݭ��� ���p[��(����G��2���B���9'q�tյ��*�����yYjP)^��W���z�Ԧ���=���ɫ�W�8N�(]�Mcz����p���匿c�06�%��Y>�/��R��v����<o�b5��:���UY>��ʋ鱗+�1�U�����O(�I0+Z�VC`���?���w�}�����~�44�Hh��� 9N���K�-Z`�Q���C��U�{��W�5^N/�U=�8��"��s���|#���Kc���c7.�\�ɵ���/M����h�ַ�0���n�_�ɷ4��HW�IFI�]kWhЭR�5(X9`Q	U_i����#yE�,���(�3�����7����YN�83<���*Y�iVa7e�����q��;�=}�r/n�ά��	:�$�9����VM秪�F'T�2��y��?�j�ܽs��/�Zd�W�(� DjAL��;"X�ᣡ8�	�[�b��#0I�Gtj�@��������h%y	wm��������-��w��{��(mO��G�}�KO��Elq�o��iz���޳{ﮪ�(^�#RB��2{��3ّĘ�ۦ1�{3ҙ
��=V^����7�B����+��A�͑���޷��C����A�dJ��S�;���z����<t�(��v�&����uI�ai����LC�4��q�w��_u��qF FB�[ġs6_UJ|�5$f���(u]��nZWN	��o�����<�7I��z~y7�OF�p�W\���@Z6�|�1].�*1�/߄V7���Q.�6�V�eN�kJ��N__|m�h�ԓl��M�,���T�����zD*�z��g���������uE+��.���C4 [6鞼�?���[�!��2f�xs�������`0桊�-���8F��Ȏ�Y�=�?\}�	����
Na����r�� �E��Pg��w��7D��->?�&���ɧ�����z�^;�H�N��siE�_;�^uj�V��}1��}�?�P��5p����\�~8�zZq�{?y�|����ԇ����gy�����?���W�Doy4�vOj�te���ј�ѫ�Ԫ�ұ�����]��d9{S�{����I|���|�<.� ��[٣7E��Å���_���t��U��b^LӃ�l���k#��smU���z�'U��J�w��ܒ_&�Uy����d�sT���֍w$���t�t��x��2���7��Ǔ֯O�hT�e����W��wqFگ"]�/8���Xޏ�<��n}�Ϋ�/t����H$��$梃S;��7�r�����=ç��u��z��p�Y+�y�_���Ut���7?R;���B?�<����x��Zp��=�,i��!a"[q�15�5mj":C�$ ?a�Ȭ��I�^�2lڢ�v�t3]$� �*䏈�s��ǉ�5Jk�pa�+�������?ګ�������0~�߹��������޵?K/�x�=���ӈK��W^��}�Ucz�^�g��w�{�����y���w��S[���{�N�<�#��;L�����d��w�o+5&��7�0��>�t���I�Vf/ϵ���a�����'�V��������LF��%��޾�{��+i=Lv���H���uN+s(@�y��ԯ���AcBH�Ii������xR1��+�Qِ��	ʰ� N@�N�'Mu��ֶ;"/K�Ә�f�6���Z���	����R�*[�|���;q��
�U(�Ӌ+�n�F5������|*⺧�A �ŗǇx��b�.��=XG�;�f�>�t����/�����o��on�	;�]#�-��l��W>�S��G��*{��h�����@V'͆�eUJ��V^���~���[��o�R��~fI�5�-r����u1�����`۾�� �s��*P���>�|V�v�g��p��ϛrE(��z���ؒK��8�����`k3�b�c����d���Gq�OB�LCh�{:�́���K��^���myW�����\]>Bj���z��Cބ���j��J?V����B�{�O�1���W:��!.�VY�)sq�ۛ�����~�R�߯z��>�/����}�p�����~�6���~ș8Q˶��%�jS3�'��Өغ�2<���,ip�Sӳ�Lޝ�3���Ԥ�n����m�H2"r.�B��m+8r�8�I���"�c����b�D�-�c �{���þKmr!��!H�=G��<�G'�&����-�M>�#��廸���I�&)�=y������ڽ�͓�����j�����_�Yp��P�	L Ʋ����Vޣ��>�t�}�~��|\͕�ا�έ�ɉ8�|�K_:|Ƨ~��-����=<��o�v��_���ĩ�ɣ�䟊��9`�p8=��,0]�eñ���{���OfӚ��L�'
���'�>���3�eH��T�%t�}/���uƤN ���J*cdӿ����B���!��$4�F-�1��oN�9yY�W��?O�D�
�+X{�L�b&�UNoT�`y����������)�P�?J�����.�����O��Qo&8�@�D#_���UP}m:<}H�K��;ʂWe��.������k������A��S�����=ï��~��>�6�ptq�[�e'��ճӣ�������&��ԫ�0 K�o����(���h�_��.�^^>2�8s�� ���( �����}��	ө�|�y�
\Y^�s?��>�ޓb9@(V���oz��7�u��}�~���=o�ɟ��:�#,.�+��ʸ6�r��v�Gjh�z՗�hl����;�����lͭ����֒��	��E䗷)��1��Y_Á)��P��z�����^��ڜ�.��?tl����:#k|o~���[��IɰC�i�(<ZA���v&z�s����$2&FGA#��3��չ����z��/��jHg�س1���_�_;�c7
�������{���a*k)S䰖<���`l��q�F%�]㣚���S6b���'h��N��ر#�w?�  H�!oT��Ґ��g�7�rg݀mo����l~%vR�:G�����[*	؀�U�9s�B��;|�w|{�Nk���?�#����	���ј���{�a��ī�+��+r<�E`�����J��^�A>���J���l�:��-��]��L��ٟ��÷��簊?�?0��/����_���b����3_��_>�������2%��0�������3)-����*}7pe�y�q(=���՜t�/����������-�Z"~���_��_���0Ҝ*��8T�ip5H��aS�{ev!���q!0������1���ܟ(\��a�;)�rP8`��X@b{�:�L-���Ib._��_��E��d$�{2�0x���}��8>�s��q�)i��HC�k%�r�,�G��޵o޷oms����^���d�_�_P�Ol�Ԇ�V�W�o�=��՗���>)�`r�]���O��=�)���\��;���%a�����;���m��.���ۯ��a����ׇ���/̱#�~�~��%Y��K��8T�B}�O�upO
��Fk�|3=�י��gsϥXC��l���a��g�<8�����m��c1���b5Qi�/���S�����-��nY�S驯�b_�3�ʋ�ȝܰ���G>�3�m.޼���� Pq'�K+@���y>[��ǜǬ�mo{[I�8����˾,��;r��㱶L�|�wf�ǿ�3dXItϘ���.�3�z]A`�
9�k���B���g��q��|���~�T$;��E9�:�����g���\}���r�9�I�w��g�D�x��v��������C�E �x�;�#Y��ַ�%R}e������P��?"�_���}o�+Fcʿ�Q����v~A��u_-�����w���Y�n�������E�F��,g�:9�J�O<�p��7���Anػ�+���iП}cL �&��}�}oM�ϼz���7g	[�2"����?�����?�;<���°�BL����W�{@�Kna�U�+�>����4����>�6��ew�ts�4�o��?���I�?���5$�+~���3�п����YHW#�82�V�Y��&Tp ����XjFk�d=�Cf:i���Dv��xu�ո�y���Y7�gk�����#Q��ﾲ˷�H��h���3U�m��#=���O�VNb6��ȍ�2	b"d5�|=�g� ��I\sX�c9~��>0��������^�ۤ��^�d\�V�)����k���M{΁����Hە���4��Q/Wt��������<�T�O��ό��[�\j�C�X;������7���R��TK�Z���.��M�W�I #^�f!��ɩf`m� �r�>M-�IO,%�'�yjT���_��+�W����K0��6Z��A%��ظ��a�GI�d\H��*��_(�6�7���&6���w����_ĕ��ѸH��Bڨ����׿\5��J��,?ݾ2�{�Ǫ�>}�'>88�@5p�^V�zW������o=����ܻ
tp���A^��J6ݜK����|G�Ͼ��/��M�U��n��v��ʍ��F�ꃦ�VWe;5�۾�j=�|������f)o:rc�{Q���~���9��Ï�~�A�B��W���~���6r��Ɋ�$�.�I"=�������3��;�DǛ/(2:@4���>$Q2�,W��BN��� 9J<ibU�D>���v"Q>4<�O�@�͒=/Ӿ�rP�#a4�=�z�S���aLi���eԔ.�FnJ\�����[܂��`^�o�G���nd��/����_4���Q�W^Ș1��).�	�|V�c�gd+|@@���o��OPʋn]jNf�o�*������/���w��� ���k}��~�Wf&pf��_~Mj��z�R���
�wW�m�{Ե������
���c�Y>�s>o�_��Ұ��ON��3ܐ&��<���{�뻇;��$q^����4|��}M�ٟ���͎\�p���1� W�Oj�?��)\�sOM�9���r:�v��ԃ�x �k�u1���R�[�,q�}(=7 u��W��v�l�a��� KE&#-x���^R2���l�^��/zQ��㮝��Ï>�ٯ����1��e/)"p��������%��}5�Q��'C��i���=WL��c�����%1������J{��r��w���QJ�!����=�V��_��Q���    IDAT��n����+τE������ַ�e��O���<��#�Z�VQV?��O{Z��Ǉ��h���=�%��ww�R�w�F��O�Hh����j��v&����e�K�6��~��_��_�l��^=V�;I���oƔ/]�bXLj���P4��zFǏ4&ox$l���o�Lͦ��i��̮K-�0��r72?��|��g�����)M��*�Uӯ���Ga9�2{���
�Dc#G��w�n�P�|K0�I�\�<z�C�4"HZX̠o���n�0��$��BL�4%+����_ؽ~y�K���I&?g]�G�!y#�������� ,@ӿ�Ù�n�����Տ�*����dS�R�)��kȮ�<x
]��wy@X����g�}�;��[�7�H�����|ӑ�[n����� ��F�������B���58e���3�4h�0Q`h�a%0�&ϟ�@���kH��	�ӳ����������wxg�"t���i9é�xb.6�c����o	i�S㔎O`�(���[�ի,_��y���z8��1������ǎ�i��/.�wI���%v	٪� �Zu���c\���m���5*�;f�����
�Or�߈�@Lg��wI1�wo�C�u�a�~_0���gc�f]�?���CA��p!'<��廢,?>�$���<Z�1�ܫ�?���V��	�������W?�_�x���w�u4=ȥa#B���MpX�63�6i~����п�|!��j�,K��6�z�k��_�Aazk�&�^�������� �ıJ/F׆K�DW�xG��l�܋#(��zF��3�$5pV��|{��\s��ݙ�����(�!�I%�
��ݥ��{3=�ƞIdȃ�MDZ����$����gϓ`��ݩ0�ެ��Z�r�ﻟ��&r �#���LcVVkdm��۠���t�X!�8��m����{-�*ǩ��6b����[���x�x�.~T�b:����H�{ۼ=ߚ�.i6�A43�:a���������O��텃��c�|��7Ǔ���G�j��kJ�+�yO5�o�U���i��L�����>b��9ٍg�k^�K�'dy�������H5(0��� [����(匟sΧa4o��l����IŏB�Uc��O0eNN��(X��ӱ�go�ƶ5���듄���|�ȯ��dN#LcQ`�ӽ�]G�g��C�F���I �2C!�OB�=�:9$� ݴ�]��U{�a�K��A5/�2��_���3�,^�^Z$�j1e��^8�'V��4����P0X����\��-�{���v�v�mW'Gj8���=�B��oP�"(�4�*�Ӆ�Ue��Ry+��wo4�3k��yz^m1Yv�������a��/��r��+�\]<w��P����ϖ�O>�\'�6�ԊW8����N���A819��ẘ���ޭ�L~��v$�AGH� ��R�0F�f�1k��vk�Al���a�و`�ࣙ0�v�M��t����2X���ЧcT^#r�F��b�eOhAtG-���J3B2����Ԣ��at'�Y�D�Y>;�n�r���j6���9R�zT��p1ug;/�>_�m�U���I���xR��Y'�k�Pꍾ�#��<�0k<�K7��TX�@���icN��վ�[Z��<&g�ங �0<p5�쵿�_+�_~�_�A��	g�c������έ<=�\��g�Q*'|�� ~��Ō�0 �M��Z���a��y����#�6��O�����D�k�P�0ĐĐ��v�&���d�1�JBZ뮚����#�H)��FD�+���a�^�RMO�>dq�ԨEy����Y뗆���̬�����c�vG]��O�!Y��zzj��"����A��N��/�y�H�yO��t*�qL(a�����x���𑴘�`� ��#�yYL�Ӡ�.x�Ȯ�c���0��?u2L�E������ޙ�	������	�ݎ/Я��o��M���]Ϥ�r��0�Rz@y1���2�3����'�����mI��4PyD�f�Y��[�0Uë�\/s�����V��R �}T�=qi���:~�x!q&-�ַ�đL�$�_J�O��v�g�T��q�Xf�G�ϓ��j0�/	����g�K��0�l'`���{C�W�1�&�WVNֽ�9�Ue*�85&�4ճ$�Z�Rm�qb�|���V�_Q	��`���J����d���f7L ~����}����`�)��1��W�8a�8aϬn�\��ܘټA5�0#��;����lcv�C�P�E]�7e}$�F����z�a �F��H5>��b�:w�lᔰ��	�C�r͘�"��N���p���Kq�:Xyj �"�`�Z0��PL¢g����e�F$�n.̡�ui� h��fU���~v�������r����R'}h���r���v+]�pVSS�1WL99�f����AV@��L�t ���c<�Y\j��z��c��`�����5k
�|k8�BzoԞ��BL�9�0;��j��Y��1&k�ڪ���Az��O;))��.D�.=8���2��`����$(ݐ	��;��&{ab�$�3��BL��w����1IO�b\j���ķd'�����N�lG�۹��!�.�A��Ԑ�2�_T8�j1@��աzb[Dx9
�}SW?,����2w�ڞb�Sz��J���tS<ƴ��k����R�t�1Q6�2��z�jĭ�fT�d[��Șj�b��"Q.��Y�:������� ���ވY�Y���F1��ҿ��b���gWwe#6SJ�cV��-d�ާ3y����%�4��[i�lX�өMD�xQ�lS�<gZ����)��E@I��*����	�>�`Mo��*wz衪�S����g>�`�������^����/|�pv�����ǆ����j��;�R���A������.��}�{����>��k��b綀��WN�>QL�LkSL����=�����}[	*s'N>V����%�1<P�r��0��l7�l��o�3�.ޓ��e&�U�H����B���>�qS&N�<=����(�����a)���n
��I)]lx%z��X�F��'Y�]]=Y�l��t���H��O���*��Zx,���3��G�v��
o������i1�q!2���EV��S�ɳo�!ܖ6 �VF�.����$kҊs�B���F���	*�S��S��J���|�5�:�8����>��컟�n�3Ir!|S��^�Χ�5�-.7%_�tV"�����|�wg����yN�>�y睵��ƛ�S#�Ǘ��*�iO{F���;�|h8P�W8o��o��z�~�^l��mӱ5&�:V���?����w?�h��OzY���0�t䆚�����\p�n8�	y����^�&��Kʅ��~)0���C~��ǆ��W�Z�3?��´��i�ǆ;�s8u�԰�/� 1�Y��-�^mƒnM2c`L�`����U1��g�v����dH�9I��$��K_2�쥟8�IV������m�҅��h�!`N����gO�4�7�J����|�/��Sgn��yW'��`
���c2�M�O9]*H/���2����.u��}D����Y\��AI
?���q#L���X]��5asۭwd��=��T���bq���RU�?�̙S��q;��p+�"�9w���$�:i���f2O��PT+xbb����n���9|�wwԧ#Uz7zV�O�M@���I��#s��2�����
ZB b#�"����b�����~��|8��L�F�=�����с�y�~�
?���E|:"�4���0�3�۲�s�*�y�`{�b�0	��g�df<KQi0���^[?Q:���_;<��G�,M��A�����
�r�b>3��L'�_L�B �:73_y{��j��ܳ`·���Uo��M��̴"��7�T������9�	s^H=��L�K�������?y���[���Yׯ!�z뭥_����5�u�u�Z5e�e�|��B��p�L5���� q�\[�0�5�'3�R_*����U��\z�'N��i�c�@���p��7�a��8Y���M�&&2�N~��O�˗	����Gؔ�z�{j���}u�C
&!I� I�id�� h3�����vt��<���ܘD���F��d�0dC`�+�8yr;�a��(}/�l��
.Fb�o�Yg����K�=�k`��w?>�|��B�z����s�f(��ԏT�ٳg�T
s�O���~�=��c�d0����Ԭ���յ0��Rl�Yf�05�y��ß��ñ>Tyr�GT���OD�&�KÝ�5[H�������^u�!%�L"Tc��v2,��m���a��c�c,�y�*377�0<����>������|K��&��L�W�w��a��2��c��58 3:����ܡ���L$��f,2Q7W�Ŭ���O��O6S�0��Ӳ˙�<�S��f����_��V��=q�^�����B����Ioq�'b��$��*L��Ku�Z�g�DT�)]1�kS=�L/�"�B�1&U�1'!쾬�DdV L�����՘�$x�Ɋ ����������X����E�5d��a
�D�+K�	����S78 �r���b�L��iې��Vd��'C^������r[�Nx��fq���A���ΕݚiV.?��psq9k #,8�	ǎ+�'�-q3)$?*��oU��.u�3p����'�����	�(��⻸,7`�&���F���1�vUN����S[f��?���/^<�>�53a�0r�~Uwڐ���|w}i��=t��0����������
!,�N<^����ʦ?�]=z$��ܼu�����~w��x]嫬�GW���S�����t�✄�{�J�3M�%	�2��0K����h��9q�������VT��M��3l�$]��f:��8�pC,� �<u���O�����	ʜ���!]cYy�Ր�"=S�����P�'X1�c�Ϥ�2HSf�}�3xNc=x�p5v3��F�iu����6���s�:��n�%>�Hp���Y��[�{�bNHH#W>:����Jo���*��2���䙛�W?+�>R�.涅���r�^�VP�� P8)֥���NLGVo?��O����Z�S�.� K7'YI)W�R&��1"�=�<�NBC�r��Cplj�lka�!T9�0�U<��}������M�THM�N8�����1��+���"�y~^�Z�"�M`�><���C�c�b۾AY�Y�M�M�I�;����&❧̩H��b-��9H�KM+c0�:�^������}	��|�����{��b4�o���LV5S���͜QC��Ou1w�̰�ṉ覎v4���{���C<���������=�2��~�a�������]����b�7Gv_<���@���j xf��G��Y�2vlf�w����^�BI�t���|����0�9�WQ�^��7{��/�[/�N�,8	]��g�6������E7�0G^���������V�X���%SFc�ѻ�DP��`^�k�>4.�����Rl��PK�OT_\��zZ	&����~G� ~���a�e�&��'��_��:j `0}�`R8kj�P=���^���翨����_��eW*+_���>�V>��\,A�(���E���ތ!�1/F孨�幩���6�s=v�ԯ��l��<kϓ4ДcH��Z�����\ a��U�<�q����O�8\s=zr��Cޯ�|d���X��u~f�>���0]�u���t*����}1E�I:�F��W��R轅|1%D����`�����.+�4�7��ߟ��%/yI�ʚ�f��^�3y������/���_�6�� 9ԃٽI�b�b����YPV�O�=O:0��l����Ņ���ȏ=�h��ʛ���{���(�U0��$�;���b��0����\$��}����V>�Y��A<�`�)1k*�L�p���5B��exzWw����m=�ͷ�:|𡇇W}ŗ-^��7V>�}񈑣�\�9�����<]s�&_,^ԁ��*e&Np)BE�DBc:8S�*ݺ�6���xf�N�j�'�"�H��$�쳚:̼�U���n!p1�w�nÌh�]#{�A�Z#�I|���_��@��w����z�ɟ�ɕO�@@�ӹ��2��ꩧ�^Μ8Y�l��d�88���f�FIKRo������E�^��G]����G�_
�F��t�r�fq���Ï{�[|²4:7fꖝ?���n����?���q%�)x�F{o$�Ñ�}�,�/Ʈk���tڢ�F�h\wá���_�=�|;��o&q�LzDuRi5���AF|{|ː*�t�1�4�F�c��b�cY�s��O����bHa.@���d��Fæ�U�W��K�U\����ڥ b4LAo�������ݧt�G�g���f��L�]�|L���e�|����<z\���`\�O~�X��&��V����Itp=�YϪ<xIH�/3Qp	w���;+ǽ�� ��]/�������T<��m���o��o��"8�f�/�@�s���7ɣ�r���{۱y/�G|���׷����;
�˼����H��pUpnց�����.%��RI�{��jW��������piĺū�@*���\'$�"q!B0;FAqUA߼��P� ��!A����xؚ/��aqC��cV�>�"6�)��\��������m��1I�$�;1KF^E5��I�ybd0��� a
���l 	�Sy��lM��D��q��b�^����|����/oD�_ǗzHיJcg�aF�wy��3���wS3��~���C��O�W�C����|�(̽g���+����NX��Q�$`#@�O�~��pU�<���:ea'�M�iѓO���p]�[�ssM�Z����R � ��š{A�{��'���Ge�w���U� 2奭HG�b�*?i<K��}^�꾥GX����퓢�NT��y'/��8|򐯺�/o�XC�W7���=�I�����m8j�>l^��Ă!O����,Nz�p ����\BY\�+��dA�^�Ա�ȇ����~�d���p�'��W/:�{0�]\�$���w�������#�F6��$��D<K����ٕl*㣒��~�n枞ܳBʙ�:x�@DBE��0�4��j��qk��@*���a'�	f�*KM�T�X\�e|�ffS>��Uq��)��y�-e�����
LZ`w/�l����IR��R�}�O�W6b�N��ʛXjvh������V6��[�:&��K>�3���w��3\��[�n�!���Jg6�@�����\z(*ޅKm���R	�0+�EP�^�p��}���7�T�h
�u�my�$wT2��+�oG�c����l�ds����Ԗ-��L�GՉ ��}7����B�]v㬅�?L%ﺙ;��A�M*kUղ�PHѢ1t�g>�9�'}�'U7D�k�dIX��b&?�c@f�)��o��o�Al��=��YX
8"�f���ַ2�M5k��;ߥ���㝠���it1V�&�|G������`$!)���Oy�]]2X�Ay���3��g�E˳M^�W���Yj �I孭���`J\��:q��W[l*�:;�L��H�����{S�ʿU��-l�4�u'ܔ)�{��N�i������|Wwxڌ��_TO���V>���]Y�X�Ѷ	���?���6�XP���~���mA-&aM�k��(��1{]�T�p�D��>*ܙC~;;�X-�t��Dب�،-z@8:,�ihn���1�]̔9	a1�[H���������Ǉ����wv�W��6-i�ک)�V�Dz!�ɓ���
�w/�Ęm9����F����KM�PW�~0%��zw.�򭺏��덾w�]́CL���1R����@wT���27��_�,��C��y���9e��Jởr��d~��ձ�%�y���3ñ��m�V0ƹ�Y�p�    IDATtq�E�[Io2��g"������DE����Z;u~�;D��C�tԃ��B_  A�tT�k�g|�gTe�O� l������&����@=���]�3�X����x��|�^��1-��@1���>M���ǤHغ`�p��>'�tZu��ީS�)���
�3��OY��{
i���k�]����MYʁg��h�SO���x�[���o��֞�C���ys�M��mo�����&��� .���{�a[Yd`������pZ��Qm=�7���X��wzo����%w��c��`�T̢p�X�Ŭ|���l;�=��k_��2O5�Dwm*�Jw�v�L��A�!D@Jy�ePF��C�b֡1'k ����-�p����7���n$g:�N� n����� b ��4&=�qkWV�	�p��y���ş�3�̅���Fm�6&�Z���@�Q�J�gp#��˦�� ~y�C��5ƄRW#�D]0��0K�C��&T����y��G8�=F���i"�L��S��z�%DF�tu�'8��5�&�¨�6N[�	q-��ؕ &���튛�U��&�o���%yL��[��$�Ǐ��-_�0U�	!��Co���AtSMvK�
	�G�����OG�4ߕԇiH̋ M�kcn��ʦ�RH�4�"*�aj�9?U'��4�λ�1R���a4V�w������\fW`x�N��d���*����3��{��Ge	��=�z�y�'��i��Q���]���=�Й<��"5�Ӱ|�HZ.z0x���3���k�N�h�<�盲HO�~����W�Hs���6�,��7X�0}`�Ѻ�wfӝ�����~��p#dv�\�6������^�Ե�eTN�rl�fT�������'Δ]���bOv�Bx1�R�H����2<�݉�*�Ņ�u�͍9�s9��>��>$5G��3a�������;O�ܔ��V�Ӹb	����|n1z�v$H�Do_�
3MD�υq�3���Ҫ��w�b�*ͬ9�}���po�b�����-/ݜ�"&e�հS�]l�N��l=B�Pl�f�Y0̠S���~�������`�Č؊:d��a2�;����0��fEL~���7���a��N�������`�.�g�ٔ�8��l��R����q�8��̩�l� ��x4n���HW{��/d�k�F������Mo��o$co��>4���?��GR����lK���L�"�H��R�)�H�npk���嬄��B�����[��i��Pҵէ�9>��8��"�쇇&^>��G�&��,�!i!���V�֟��Mri�Z&����Z�����F�)�߿�67S.��8̍�+�Q!��NV�H/_�%(�3���9�I���H(� +EF	׶\$O�ϑ,8eq�$��J�Eˋ�3�"7�v�ӳ�<;��t|];�-�8{��HJ6��V���y*`U��R��A*���3���
|�j����r���,�=w}cex�3��_V�\<W�� y+S��b�V�=:}t�>&��=�sa�H��������)K�Ƽ��v�ܩ�jȔ��JJ��e*����u.��_V@�id��h&W=��Ne@I��c���9����@ʣ�{��ѹ�{��H������f�z(��?H�?\/W�R9KU��S� �!�F���=�����ѧ���Q7���m���b���_�j�H%�Ę&u� f)��u��?�Aˁ}\U�{�Y�ɔ�N��EB��J��H-Ʀ�|�me�Y[��1GE���b�\٬|''V�^�g0�6Mn�Xوq!V��Y�Y*@V������]ԣZd�!n�����:�;��f���CK�5���~6W�~���b����9�6��x.���d��?�W�7�t} T7�=Aؼ���Yw&�s`x��4��e�赳�fz���Y����l|y���ИW��pg�w>4�K���2� wzo���=�3LM-��9�{���|�~=�v2��O��������CZ����a�ލ ��
���5���g4NZ�	<��q���.w������/�/rH��u��Ȉ�F�=Db|2�x�U�w��rq1��L��ed��^��Ft&D��K.�dƴI��ߎ��3�E�u���I��ﺷ�˂i
��)y$ݷ�51���
�z�ɤ�SҒi�nX����ұ��xs<�߅0��ӏş�Ψ"���I`��
���G������Q� v/0��RlõΞS�-&̪&��=qӊf'k��ѧ�����Q�Dz�Y"øi:��	�R�4�������۲��7.~YH��x������O�F!��=��͹���^?sOd,c"�*љ
��r6���~����mk��l}{`1�	�=xv2Q>:�=�����k2-�:���0� #(_Pfop���HI��@���4���a��mne����t��?�>s����ax�;ޞn�^})=J,9�g7���3y�wbVz�K��P����I�+G�ə0VtPD�@��&]0\5�FOc�ы��@=㖭����s�3֘�}���X�Ƕ����$��]	zШ�a\� �@Ofܠ+tf�X����gQ�,�)t��{"���3�bf��H���8r|������S��o"�e	�����L&C��/�˧��؊��L�;s�ԥv�M���wT_��9�+@()i� P�u�C�F] ��j����./>0�Kr4>�����~c|��L�o�?��h���6<r��4��OR�Z�Vq倥36��,
�6XL����</^��i�s��������E%��r�+�gx��o�r�����F;YW9��#�2��������i&:����$sr˗����0�D5x�4+�2pԣY�y˭7�w�T����ca�>g�!��,ڥ����o�:�K��q�ʇ�Vf�4F���Zޙ�G?��;�Q�0	�{�k�Yaz�jzF��O�e8�	����vr�S�>;���s��إ3�1�Mdq���[����h	�R%m���ۓί'�O�/�G�u>�#��ѹ�����~t8�K��f�T'���R�ŀK٤e%��\*�E��]�����GO�S�}0*E���d͆9����{�D������".y"b�ЧtK�tx�@��I
#�6�� ��/=��lu��t���><��E�=~��񙅽s+K7<����qx�����v��n�	j{`k�o���������6]c���$4;�r16ɮ�!�3V/�������v����h3�5�Lfm�Dc��>�y�3��{�}-�w�+�̰C�97U�0N��a[ωR��=��F��e�͑M�~�'~������Xh���SqZ�f�'��>t��`9��U֨g�	�24,o���ն�����R5yAR}�ę6��-}#�/�~��X��0\�Zd�>�c+N�Y�ވ�~$��	Y�#$�hV�<ЛuM�#=�h[Ic�IȽ+�Ҟ��g�$u�R������p����|��F�R7Ds���Ƞ��T����y&a���t�`y����3x�i�$Ji
m�Ù����Φ+����ٽ3{�9wr���S�-��4��7�r��I򪃺��#r1Ts��}ߌz��7����1��O8�RQi�nW����2���'>e�=)n+����'����ު{I���Pp/�ш0�F�7{���ѯ2��Vgz3�S!�3مц�`)�V���r���s��Cs1�M�ʼ�������G���<s�Ԥ��3��6����#ێ���d��YK�Ӷԁ>p7c�ë�N�����c�{����f�">�����̗��\->�U��!�$�.2��
Bd���䱱�NY����}�Y�[����k'O��̆/��A{h�-R3�ɟoFR6��K��*�_��e��7�DX�Wc��㫑�����Z]����H�Ŵq!��}ss�1�/�LxaJ̠q�I��^���������~�NoC�JRS�����=9*�9�l,�ؿϞ9�squ*�'�28���icnj���ō�?p�o}k&B�H8���p15�Lo�5&7���z"�z�7���F�+��YF��4�e��2p�{ە��?�����K۟��>�'N<~8{�L�p�fj���n�p���Bή�>���GP4̠9��Wd�2���O��g`xE�k��f�9gH�j�1� yl��mE�9���G�sf4"_�����k���Z��	 a��)h�����	�����%�r�Y��)*jCt�c��0�!�gG?/�-,��ܾ�ӳ7�tˑ�CSQO�]f<HBL���<I�����2#���ZE�q6���w��$�%P��e	J_��'Oon�.-�lLL�Lf����ٹ��{������x��K*v\����t�Hs�2i�z�Dj�SzyI�H'�6`�7ͼ)�9wv}n{ϙ�3�1�������'w�N�n�D�����֞L�M��H
k�;�'���C���춘C�G*�l7���>&���+��]��̧�΅�&�{�o,��ؙ�Iٿmfyssgn+�O�XTM��0&-���d�2:���@�����Yi�.i6ih`�j�>뛗67���OrOl���g��������z�0MB��*u�,��X0�k�tS*�XEUx2�h]8��mtm�<4����,q#߶S�����w��C�fl�v�"1�.E�f�)/���P��U.�8A
e��6��t��0���T~f�2�����p�m���^��mN�m�Y?������d�:рL�'�1S�HP'x���`���tpfѭt�'�4L���0?+�U"xY�Z߼0�x`}'{O�]�ܘ�[����{�칋w�F߿�HA��z���5��&s0�F�lF
ܙ����D��M=���5�g;��&h+Ri���Vv��$��wi�dTǙ����'�/\���[/��l��,]�w��W�^+p���|VU�����1��3���qqq��㦓S�B���$�'����8����!�y�����`y|C�J���&D�����6��:S�p���M�ܺ���?k�#7]���_��޳y��O;��Ox~I|]�AZ�!䍉����m��	�����nNC@t0�8q���F3"�b��{��ژ|���΃�k;��V'Xߞ|8��^HCٱ�K��h�=�<�ԙ�;��x,��ݲ�l�A=~_��QA6�m��>�|~����2�����(��֧c�����/�용��sv�
>���-Ѕ<���ԡ�Ϣ>.?���]:��V�������KS{�]�
+��{��ت�9(K|�k�)�\Fw�v�#�\�b`h�Z9�H��W�6�� ���������}��-��0�}�5�K���!� ���������`Ez��fPi^����)�߰6�pxmz����ҁ�#�=���LMo����̜��B"�� {|L�!)��HF��b�R>�$���\�'\^�=��6������k'�6���{b~~��lTp`F�s�i7���z����I���3��&�U����yHc��u�ңŤ~a��օ����m=�j<x!������޽ϲM[��V�0S�f�+�1X���%e4����ϺJ�Jo��?*�Y:LP�� ���,e��g�7^��l"�ށr#s��[ۓ���Μ���3�͚�� Rwu�wM��'p"�$*A���i&-�E�d���I=��'��\��/�NI `p��жPݲ����&4$v�7�}]%�?��U$��p�\Xv>�=��V���,�GzڰᔣA�À���ș�C4pv&��Q������յp���nz�͜��_�ޞ٘��<�g��b�&Y�fg�lӋ�����5fV6GT0�jp5PJ#�p�+���tM����9Vzeckw{*:mN$Y���z$��F�S�/�L�xF\f4S�2<c� ��Z(�,G|��l��	&[����z����<�F m��~��]nw6�?���/��5җ�VT#�*���p��P�{�\�C;0g�"O�k� �5�c��+�.�6��[�%�I;Ƃ�w�=�xf����uUwC�4q\uO2sy�wn��n����͘��Pj6JyVi�>��\V��:5�!F!:� ��w��t�9�C�Mg �j�L�ą�.]��{�衻�3K�w&��9usb{����|���}WO�>���ѣk$����:B���O�~�zf�^����2�8�0O]#ť�PrIqM�]�ڝ�>�y��I[�]�!�s;��/d�l�`^j�C9�u�QM��P���x�iO�k��o��{�ynImh��ɴ�)���{k	O����}γm|��ęǟ����s��#/\�p��˧�w��cύJ��^�o�:���4��^������z `�<��5��iqa�̥���q'��AO��Z�鹷����_����s�V^F�|���F��ٔU���~�g�$�V����񇫲��K�]��m����;9�";�nf�y��w�Ο={0�*�:}j>��5�������)�H��#S�����a��k����،����F��_�ar��-7�\�V��.̬onN���w{hyl����e�S�졝��ǚ2��w�k.<��&m����w�1r]�}�;w��{���7)R�$S�]S�,)N�q�T�0M�p[@MӨ�?-�4(� h�(��H[5i���Ӱv�(�r�Rd�R���II+r�%�=�;s���s�^�bH�"��V�^i8����������A��kQf�@|6�駟NLN�H���|����f�TX|Y��<s]ŚpŶ�:�-j���R�r��6�7��di���ā��X#z�R�R�<Qh&����hK	f��{����}��g�]�w�L�<��(+�1Y����Ɓl~�c�-{����6�0a�z�x���M�5k���$"�S��㮻�2 ���W�b�
p����#��J8lZ�	�?R��[��`M!{43x�?w��333�v*[�����Lk
JP�e�f$3.�� �۶�+�T}�≉Y&+*A�e�-*�yQ1?=s�Tz���>2L1u�������u�ًsBL�m�`mRb�ǶL�vY���2�9dâ�s�,�����%m�R��._�|��E�2�׼��{�'ƚ��.z��۽�C�VUe��m��s���FǶ����d��������Ǹ�ey�Ȫ�Jg�)��#O��_K��ֱl��N��.�:h�����.-�	{0~ Š�r�};�O�.�-"�^��蔇�ؘ�V{ep��6Zu�-	��	������tqr����?��W��+ SX�_�N�W�.'��8pŲ�d�.����ժ����x��iYX$Fh�iwmɲ�Rc _��2
��z��:l�h]Qq��H-5ț�\v�=?��x饗_���6�7�F���o��9�%���w��O��jd/�l�8}��#�ꝼ��٩;v�=}���f�C����"W�쌡ZP3dbX�7*Vν8���[��8�de�:yR ��w���I�ڔN�.��fd�IcWd~� ��S���g����QˊmB@�����|�TP�P��*�R�R��vT��qT|'_�9�e��G����<s��lO�K�U�v���Vl��^����?��ta�B�M��{`!��}(7A�
C���(�j�mݚ�0}:�Ƨ�)�Zd�K�ۍv�z=){��gX:mUJ���7ҟ�X��X/���Û��2���ވ�;�i�-�	����+`	D�g��R��'�k�&��ʘ��X_�M2��@Q�e���*�,��X�d��̅}A��r���7ҹ�����z�����}�*�����?���c�^�3&��xO��.,�*��v�#�`�>\D�  �l�Vm(�� ��P�h[����/��WYJ$��l��BJY�8�@ 2?��(�  @f����I���Hjm�<��c^��.y���pə�T/m��=��� "��X[Pt�X�i�)Bn�FQ
�����AQ�oY#�g>��9�W�YW����K�)9dp�P,�N6����;�n��Gg���Q��    IDAT�JF��ܸ"d��������|簢7˦�{�>�U�wH���Fkc��9�C��_d�����p{�7����E��r9������l�zǏ�,�?�䟵Bnco����{�wpq�U� �H��2?iU������w ,@ @E��+5a������}�8wN�r�8 @3��4����b��k��`L�� �g��Ŧ�)<�Hy��/�ӣ���G�w����.^��k�Zbt �k5Ŗ6��6D\�ܓ{�"K���8
�N�I�p@0� ��.s�C��4�N�h��rgK)i�L��Rٿ��=��xr�9�֥�Sw%J��c۶ٱ�b�8�I'�6Wl;۶;�����~é˺����c��f<����p�+Nx�
m�ѽ����(�6�Qz=��^\(DE�$�(�EB�;hL d}~��o:�x�_�X��������`��`3�O����6�H���f�k�3s�;�p)��i�{��#+��t��9Nw���YQ9H��v�J[� H��}3#J�󹴘�0to�$H^غuQ���6Z8d�����`�Lt��{*T��te�˱��	�}zuzЛh�N�y�<!��m&[���A���J�%�&��
�	a]��.M�#;LD�~^�]�=�y�jZ�lo��쩩����cJ���M�_%��x���ux��P������a��"�p��T=�(wϤ�n~=i�u�`u�`�NJ��/
��؁[�x��$�}�aa;yU��Rb��5����9Am�{]��Sf{]tI�b�� �{����ų�����$^_yC���f��UC���2�������:j��M�@Mp���̄�rɍ$9�IQ��xrp���tUP��G�PTU�VF�'��r��d(�!�p`�q�2bH�9CV�!x�.���Z$�AA1����L*�<(|Zb�>�)�X���:�F���җW�*�.��WBW� n�ƹ�7Kg�׆C��A�%X� �p7ZLL�Ʋ.�97jz6mjdit҆��u�����n~`~�P�������Р�g=O�p� }�3�ub��#��m�1�,x�M)��M��
�b���1y�
ղI�G7�L��.\�f3���SNJw�s#%��2o.��P���^��1P	�l�֩���Y�(�^w7�#�֕F$�_ή$N��{�R�.�T�J̠I;�x��y�եlſ9�5�j�������;����0�%B�zh��f����|�K�7M��jH6Y�Y"�XG�#ѹ?�ތy��D�
�e�k�����S�A4�J�)BeQf��z�!����������4�1X�کzB�g��\����-d��a	H�G�@�8u;������OHi<G���B�?V����6��D/GQ%|�	�*]N��P,j!�D��f��/r�1�鹚�;$�aa�nا��� ���t�C�����<@��a� ���ǔ�����D�xvv��K�b�����>��
�\-��4\��5������ {C�!�D�Q=B�W	�T:2QD��o����o�[O=�({+ǲ��k�~.�x�ƣ~����f��V2�`@��7�l��%������s(��z���n�.0�ٝ<�+��״�=`\��W�57?����%�e�l4S���~0"��ZX̜77F >��BOb.75���]��{���T��~UhVFq�d�R t֑�)�*3��c�U��0��uQdE���1��ڵ/�C� �IU#�gg*A#��K�� �-?V�L�&�5�"�2P�D��X˟6u��.s^�"5\[شS~���_���Rb���,H�fT,�`���!�x�O3Iw����Gr6�3$8|��D������`�!�N̏�(�������n6{2���J���!5S!NOh�Ta-��o����u�������
��[X��?۸�~啖 �k�[2i<P�̂V��<G��K��É5���FHǲ>&Q���u0�G�BE���X��Ua�f5��#|������}��Pa� �n�}�/�u|�2��[\t��O9&O&�+Lhd���rH��\���'�AX���n�k�5ĆB���g2M�[~� �a�qy��.c�����A g���������̉q��^?	�.oYBe#�O^0��_8�m7ܗ��ۦ���K53-^2�`��$1�M���M�w��\ψ����qect�䝤�i��}۳�@��r��ي��c/��C�/���o���n��5�\hТm8C��A&2i���tEi"���ʠ%���>��b��~6H�`@����.y�ة�d�n�<B{�攊9��Hb�@iS��C)�l���R���Ur����a�{B�ru�����K�H�0�*띃;<���۩���K�o�6َa�8�I�[����/����y����B���y;����QOM�t8�i��/I?k6�K�BXb�$Q�զ����tb�
]
�)���Z3>8�6�o�aV/�Ŋf���2kB�Æ�c��k|��մ,ސwR��$
���<�l���M^���cS��)�t�㎛g.�!D��o4�-m�%�!�d˃v0v�X�v},��1H��1!1uN{���>G�tz|Zp��<4�ۤ�t˞h�(�;�J��P�&>�F���1��m4�$l��2M�%�)��*J���\�&^˱��*Tk
"&Eޙ%L���u`z�;j�����	��SFQ��ˌ=XK�b��������2XM�a���$5!�jd!�Y��0	�jޓ���>�������J��W��;���7TD7����!���������P.��f���T�(ϷE}��t^�>C�����zG�pȭ���z��/�_4\s�R�hqD�,���A�ɞ�(���-뙨�����0�0&e�2���a�P��Ź*�dQJfy����_
z{�)�z) ���=V�+���U�Q(��Tsّ=\����ƂsLP� ��%�Bq't�Y���|�q���6��|���o2�.l ��ńQ��V���`��޳"3:�p�m�W�m��%_h�x�����xB�H}�ėT)`��r�2��wD��a�5z-��W����-��mG��YM5*���Gbd�zA�����JU]���C�c7����;ClXV��͎��6_�+�n��[�A��l涡$mh��6e�v�|*,��::��\��`+�|[��R����:d��Tn8�"�?B�#SddZA�^A*�( Xp��rQEv`���5�2 dBt��"�w�.:b�8(#�m/8�E�
M�H#G����I���*�b�� �(�^nͭ/-�(����yR	 ?�yҝ>��Q?�w����B�I187:�e�>���mE3 S Z��k K�2`��k��p�akBI��1�k����EVmO�\#gO�/��83��͇�a���m8I�y�̔�.���Ի�'�d����8��5̣�0S�ծ�������Ξ�Dz��v����ʽ�	Kus+�Aq�'',�Jbp\!e���i�W^J��(��ӦI�ע�F��4��9+��F
aO�jQ7��W!��:�yf�$i�S�πQ��2�Y��hk���U�QY��A�����6[y-����0Y�^ngK��<�G�+
+%N�a/�w�)O����fՂ�L��*����G��>%)>�V�ƆjFm�o@���˱��'�j�є�t8������A�z���]�-q�L*Ng$���@J���y�3-���l��pD�e������Q��CiӲ�C�9�W`'��l���y�-r�����2hEa ��|��6v|�S��tU�-���uܢ���v�U9��H�hP�7�4B��1t�(̈`��.�I>���ݶ5�x�2�w�ni�<��`T�vғE�TSi'�;�2��1r���uS�S\�.r4�R�~��+GA2����@����ܽ�2`�����v�R��'T6�β�[�:⻪�x��BN*@g��Q�|:���Cd$�w#l�zC��n�������Ae��D��(����$b����	�&5��*ϋ[-&CK�W^%Ï4�-�a�0�^��`���d (�MON�;�n��6���ޯk�Φ�U^C@��q��2s�2��7s�;'�#֒�܂���|��|đ����ոu���u�Xb��i�+}]e�=B�Ș7�H�)|���*���S��=�oz��~rdr��kkUo���TJ����T_�1�d��M5�Ũ��ͷ���$�`ձNg��xz��!p��U��,�Q�v^Fr=Re�%-��G�]Z��/kguX����=��'�����e��U��9y��u�)���	pQ�Z��L�0��tt=lo$�[�ʳ�;����`=l=���f�jX�aOHՇϓ"Bb�z���w�[R~3}'�NvL^QjMf��lD�Ɗ
��Ϣ��r�4�i��}�d�`�r��~a��U��)��V9�i�qy�5�R=R�+q�ɻ�ʹߠaW�)̙Ħ�{�W�H���	���\q�3�K��~n�E��-2����:[�H_1Dוt����������"�ܥC�ʪ�[���.H;��x͵���$�����;d3��u'�rhA�;+mwtO9Kj�F#_�b'�/�dN��X�m.JK�B�Ѧ�[�]]qM����]�1��̷���8*����oᯀ��7���lT%>	��1m���V�%��y�&������"m<>ː�Ȕ�!~�ȷ=�����+��
w�D�����KZ����6l@�F&%�4��N�J���T��b?��ߏ���Z�J;�wۢg�+�D�7�U�%BN�7hg"�и�իfXݲ�����x�EC+�}����sK��(S��N?���߽�p
+��%�x߰��ˇ>I���Ŭ�΋GE���{y�.�'�'����v��g;����R~-�9�Ju���@ֈG�&��] ��q�I�[���Pǡՙ%t��j�0�'n�W�cK}U�.�06�PwT�ڽky�5�O�+^��TMϖ�Ï^w�Nl@�ɾ^�j?����<Q����*�8Sã���~��d��c��;��M�������G5����r�p�ͬ}��~�~�Ԟ�z����3e�spF�Jmz����')בd�Zʒ�@��Ƌ�s�d:!�/��5�}��g����nvH������;�	�n
9����e��bڴ����#M6(a��K�F��{BJ"������T����bn0���a�[�M�仝���f\eemI��K��p� ��Q �³P-BKfL�B	Zÿ ٲ���8;�]2�m;W��n\K�RQY_�R"�p�Jy�w5��(���F�+WO|�5\r��1���l�E�Y2���^܇�`�F��ʠ2�:a�/��jR��m�T-�cV�(�@�Ռ�s�������f�C�_�"-�a���.������J�'�Q�MԴf�<hPS �W�P�ǧ���O��v�^}���J;.-�>��G�y���Y�H�{��#o��3�D��ɫة̫F�6)��$����*�vuT��j����5$f�5C33�&;󚙝�)R~HA!�'cf0I˨�J�ȔT�����v�o���x �@�YHa��f����.�O������k���<���L�,N��l��lI���j�>l��*���.���	�� ����0��Ի����C�6:��ki>�"��ע�[cCM0Aň�6�`�,��Mm��D�dx�K$M��&d�*E�w]K�K޹"yL��5n[ʌ��A6����+�� P���-�q�6h���4�I��ج5�'�=�&@o�U��y��DLB������;��:o7m�����o~�F�C�,�,�B
>ྌ����,�%al�e�����r��څ��?#考̯�=Ws����d����%�BO�_�OM��ë���K��6�����5兓�$�Y��_�c���;S2Ȱ4�7�s�/ȣ���IS���dx/d���v�H��R�H�F^���0V��ȏ�w`M����cF�`Y�C��\n>y����>j�,¼��8X4�QE�Cĥ8֛H;WZ	?I!@~x�8��F\�\M]u��`]T�o;P:�0��yE�d���|rĘ�� ��_��]40]\���.�ktO1,��, ����k/P1@�m��:�K�`
Ҁ��B��
M��b3|�v��,���΋���4�D!��F!|����6�pza\�%E���l�i�$U8D�Kϥ*���<d��Ҩ���nD-aRwE�.7aƏp�����{Z~8P_�ľ��N���B�b��品�B���a���L���ז�(�s-n�aK`��B���8j<E��Z���בJ	������	�%��﭂U�u�<�|?�bz�#��v�?>r����MA���[~;�K�
�m�p��3a�k�̬*6���l�oJW�n���=:;Ҵ�p�Hb�5�kw3?�U���ዳ�$��7�M�j'�q���vȚ��Ӧ�#Zz3>�L���$
��
�[��&7��E$��鐺ο�1����̠��b�����]\��'Us��/�ش3�DM���4�_m�M1��*� Qw~g����n{��ɪ�y���Ǚ��u�L�҄ȣ�G��Sn,5ÚX�s�_�r�dbmӗ:�x�6������'~+����Г���LU�.]�{Ԉ����h����j@����'�.y��x~�	_����MAsñ�6�<�o.�??+���Z� l����l/��R 
_�1.��x��ݤ��bVM,��Ҧ�} {�yi����+w-J:��'ko�|��#i,�j�8���qfhn��h�ٓ�Ԭ�{�a@B� �F�e
6Y Y��̷W�^��~�R3��St�M�Ɇ	z}�jw�aG[	_0+O����@0I��ק��Co-��X$ĵó�G�������?���d�"5�R�3�1�����ӑ�@��Y(��j�'4��	����@3(^bܕt��'qC��K�c�EI�Fn�����q;t��J(�t��N�ǭAO�$��JRO��'<^�!mXL����q�e���(�Q*�]�1��tC)�{QY[��y�M�/9�|*�t�QF����'��!fl�VK�zS�'�fE^�)(-�S*���q{H��`i��=�e&��֙I��l2q�zT5!���.l���@�	��޻n��&�O��1$�[z��=h|`̒��n�%�����7�,o�:V�ыB�
լA�`�aW=AZ�$���X���B���=`���F㚜Z	��T�i4�:vX'���!�R
����<;"�_�+n}�a��AE ��5��t?D��5��4'\��K3ɋ�M�a���y4O d���J��j��$nǌD�g�E��)��"�
.i��1��ޟ�Y(\����I�R����v�a�˞���x��TΥ&��`��
7w�g��-���y]h��1;�p���F���\K~���&(U&�<ᴤ����\���C�Hװ���4�	��d�Ȅ'����U���*�]�`j�
l������5��IhX��G/܄r�7>������Aoul�v�3��<�% � �:j�:����F5Kq)Bsc
zbڤ_���5ɗ� Ե0Y>��)�T�<P��gX��;��0K`2�]�����!��:��7A����`�,Y�A=���W"nC'53��,{�Ȓ�lD�F� Ib<OHA��tk����pܪ�wL����:�k����a4�K�`I�i]���v����E�'�Ze�@]�V9=�����dzB�H���g.�B��S��QU�+��Y9�9������Y�NR��t)=�C��
1�$�@6���/f�&hݼ� �̻C_�`mȏ�|�}�+��j
�d��&&~��V�]���]�/s6�S�f�<K�$s��Uڲ��sJ���0���C�P��̞J��|��2)�y u}s܀S����c�X܅G_}���O���y�<Q!��,-��?bgo��Y;������ []�gw����0�tĴ���Z�d�d�O�O��uQC/8�՛MN~���S����QW�X"�D�'��	ٵ.9���%��Xs�����/�Nw]�L��n����my���v�;dCF��C�M�1X�	%8�}�*&L��7�g �4�4�Yc�b�J�8�����^f&�vz��>�4�(��İ�|�	�@���Ƭ[�2�.�9��/�<��*n.���f��%Tg{8��I��.��D�c!�A�PRM��j�<�T�_�A��fG��U�*T�;l -�/-��*k��K9P�����^��j`*b��iv��IbAr*��y>aƘ�
5+� �sW��6W��	�7���^?�I/���}"ژ��.V|<:!+7.���r���^��Rk��j�02F?0���&��*�1�5�\&]]�+�|�' �\}^"\���C����
��oҚp"ꀆ`�K�(�7%O�a��l�����հ>64A��&��l��ee9q�G^���W��;�us?l�ɥ��1;-,S<���)���A���z���s:�f�1��?G� zd�O��6Ć4��zֽh���a0URVn6�И2�9��_��{)R,f�e=l�/���#����ل�����ʊvȂm��Ts�=Oz��B
���Ȑl�P�,���*��,DN*ZU5Q��>�:bXj�e��:O6O���
�|�J�6 L�,أ���GkϾZ�5�^\س��j�xi4x�aA>�T�zE��)6�&������%u��oy߽�ч������wF�K~�:���}
��[��D8��7��v/������U���L�t1�3�t�KT*�.\[C5�7�g��f�:�f�-@b�k�E`A�*�sd��o��%]J"���z(���Y��+0�w?��L}�7N�����x��GI�t��^�����Xmb���	qw�� 8-�9��1��j�����e�m��xUM&?2��1�⠋Xo���LPZ���C#o4Su�Ip�?u�~mg4�qb,..�9ΗKսi�XU��7⯢xU�ē�l`�3T계�����Z��~���i'�|P�T�+j׮�c	F��u��f�4�h0�X�eb���5����3�����4_��ӵ%�\bg\�� w=g�$�������TVR���8P"��䞂,�����c�83��qU��S���PC6�2<^8�{�6�Z-��y쿦ȋ�P���1+V/P�:�}�s�������,$��TA����Ocg��s\�=��� 6H�2�E{�)S$Em�D�k2�MeY=6�Ϩ��E=r������������	���
��	AG���HF>Ӵz�u^X[ȟ:k�.:aybl�voΖ�eB�E�_�z1�(�߾iB�O�@��QCq��V�L`���rD-E�b�r[�7�t���;�ۈ�^����?��K�n&:M��� HB�-�cқ;6^�6��J�̵x�����#�,�?��?gHy��'7�c|�>X�t��6�6Vr�.��9ӊ�Fvv�ˑ��L��6&����?��s�RJ7�H��J��b@�Lqf({��֨}Z�����{�@`Q�u�)��y(#A�n�����6��1�ы}cd	�!�	\]?�ǹ���'� -'��G�j�}DpM��P3ETw���x������^}�%$
J��7q�{6jQ/�b/'O��G��3֖X�꽟�����=A�j�b�! ~+�>t�
��=��l�@�`����Z��[�
3����=��4%��B>�C�C�#��Ҋc�S����э����l�*
�%��iUHu�3Z�#�7b�G�f��~��~1iA>���f"{9����V�톼o��5����>:�y)),LI����CG�֎���8�f1OO���m�&�7��G����	r���c�9�B�A�CО��w&|i񢒹ʹ��������ñ��i�闱P�d���P2h#���|�V,)��[3�����@a�2�)�������h���Â�<��zD(��D���̐H�F�X���Ԝy�T֠ՇprЎ�.��@:D��L���'g��mv����qanv��}�����
�F�^�fRi�d�\lxi1��P��+�| +�u�j��s��o��kQ��V�fR��Tjxim����f�q�&^�f� �B�JA�
�&�@��پ��ր�J��#"� (��"� �;�<��X` �؉0p�?d*@�&�LP��c�G�F1ϒ��N�i� ~���^J���n��:%�U��%o%��h�;x˔]:,g{�H �P!(�^��H
�?x���y�#%[�`�/��#�?aWuI�UY��w�͐�+BUg��TJ$,��I�ߌ�Ҋ>l�T5�C�V!\��<�z!�iw9U��/"�?�	��#��$��aK��1��4 }
�$g�۱g&�g2��B���V�"��)��j���W`X��`� ��c�$�t����I2��	�W���=�h+�41 ͹�S��B�v��A�!GeM?�s�Z�k�����Y�8�T�X=VB��9�d@�$�ԾLFυ\ycei*
^��Llbߴ�\�B/�a�5f�W�0ر�1dwi������/'�9����9��cn��%zR;M�΅���1o��i���K�XI�+25����6�Ae3V�g麕I��F;��Ѳ��J_����0�j�����5��ܺ�d;��j�`@k2	��`�֚)z����k�4�C̓T)�a30ǔT����~A�;ӵ���uϋ���Ș-|���:'{��]c7����*b����`?M*��c����9�j�w���]�B���=S�����VϱA�.4���?2�	�������2�GU��/�Y�D_g����K^7N�OO��'GQ��a��`c#��b������Z�g�l躚G�ٚeT�O?$H��f��<��GY���=����74�ۤ"��
��@��y�3Sה��q}5�[l5�K�6!j��=�����o�t��*���f;ZV9C��/���S
,�+ #�Lqc��F Y/أ�A�c̀�Z�У�n�ov�*W�El(�01�8��6� �;���l�
�ҋ*�uq��6�8Q�1a�ID��/���{c�$T7�'���0|���{@��D�0�䰉{��,�1pp�I*R�H�f�ş#�x9Y�nujab�)����6��ā{ c��_}	SR�b��Ճ ��}'�x%�H����y"���h��~��-�ZS�&�p!� !V��u�j��:�bK�*���y�7"U
5�D��}�F!��u��Z�*_mN�Jq�ke�\����|�Ċx��W����X���#	&��L�$w֩~<N��\���GL_�sZ���ǧ�s�*R�\��Ъ�e�*��:��"���Ֆt��0�;N�m!3I�j?@?v�P�H:~DK���"A���K���o�Am\���%u�j��\ދ��3�}��dq�W�U�a���X���rz~��c̠Z%�փ��i��pg�E�_0%�\p���X;ђ�.	ѱ!6�̄oɁ���~�F;0��{�D�"<�y;N�a�hF��#��}A���Ұ���r��`�ڞR���F���JǬ_�c?��'r���k�oh��`�K��델�}*�E�=��ᶨ1���|�*�iTn���$���x��#�m�������aǎ|��FH��$+�sQ3e�dХ�\���IѲ1"�?>��u)����Ĵ�6)/X 3�:���$΀򯻣����� ���8̫���N(�P��V��v����r�%�K[�m)K��b��������R �����_��������:.BmɎ��θ���i�-�y@��W�s!�7��ƀ��A5ȸݎ̙�ń�hb�4��9��4J�/,�y����-�y��z���kh��$
.��iZ�)�h�pX�5vNpV��G���x0[��7�tVj��D����/I�3�. �7H(}ͼ	,j����hx�q��OK}| #�\�l}��^�y�&G��?,�W�Sn��TU�g��	%B`���Z`��c���]|�1+C��3�8r�>iW�)=���a�?U��׉YT�r,�q1��č�k$�4�t�����ӣ���
o-�W+Q�ԉ����*C��z��&�7�qq�c���T`e�4,��zX�8������	<��\H}�7���d������0}U�&dE�����-FG	F�˩�����+�F��ؖ5:����	�����l^��NT  ��T�,cHzs��7Ե�40G�d_~�@��^�_�<��3S� �c�l D����ȹ����5om�G8x���4�� 6'��֒E��!�Ú�����Ϥ����r��'H�T�z�`5�D�?�#�S��%�U!�&%ww8�<����O������ѐDN�:��H3cd���|�&;�����C��v�Q	V��Dtl�qTd��bw�e]I���E�^�)�!Τ���.�b	��2�RҜm�r�~V���y�u��/�Ou�l,�;&|8���Ο5Rk��1tkΛ�p�*6@ƫ��y\L*��*i�%�;��������Mk��
͚dnï9im�(D4b���n[�9?W7.P��7��6��Nu% 0�G��WT'|
��p�#MW��*��X�4�BS񈉕�v:tF,���Tx#i���>�H_O��K��(�~U��g����##�a��l?�� e�g��u�y����)4�H�^��h������3NU; \��
��l��:y�D�`�����unlc���4��F�"�:Gխ��^[,��;L���(V�'1��W{_O��$���m��i�e��Z�m����Wߺ���j�L]�u+�Ꙩ��a��sZ&<��G8�6���E��?�>�;m���X�P��9�Jq��W����bH�y��HW��~�u���B^�M$I��L9LLUh�jQ������%�Z��@�/��&�[����=Su9(�A��D��q���v˩� R*��2�0`}"��V��n[w�b�i���躞�%&������<�����Ƒ��%:�OE�S�y_��|?G��{�(�ԦO¿�g�1�y��b�TIA sú�i�t\s�J�Ū¯�j�����?}C}��ǚ�}t�gÂO�un�4.M�% X�_����?�����u�2fD���LSg�8��\��.2���y�T����s�R����a����̌��/F�;3�7�Ѹ+{���#]�۶y�U!g�;�f��.�ѲK�@��[�0��H���^^>�%Ha�^��.�Y��r:�i�|b��t�ۮ�M��me��M�T�w5�����G�5��T���Ξ?���ݮ��n�9�"�}��[̑r�+c2�4��t������R�ǽUi)��&����?.�q+}����p��/l�LA��]��F��u�_k^��U�B��a��\�G{�xw���l�}�{���ZFj>j�VH�W8��P?�F������o���k9�Npg;+�ʉ�&o�Y~N�]pn|i���*�}���Q7/u����s���| �B���.�Y掏5����x55���_�x�� S|G܅ʶ�R14�ߣ�'�ܸ��۽��n��'�_����:�$��5u�(@H-7�OQϤ���[�z�7��GR/�80ʿ����qp�?ӈ;�g�����rz�P�ޖ����y2�K{�oVo]&������s��o�w�YQ�bԥhG�K���K1�܏'��s����^�-�"�4�.^�~̫}��Rw�u� �T =����b����|w�1�򫌻��[�:�)l�ޤ7^�.�����
曮:.֭m�g�5m(�� 1�Q��ۜ:�6�>#{}�n�I=ob/��/�'��Jo@SFn�-���5��Z�ٺ��J�K���6����>�ﻛ%�E�,�(��fA����Z��˨����v��J����MMmE�X]���˶{��+�e,�g���%Zl��Y�4�N�G����x_&ۗ��vU��q���y%_ga�����\��c��lO�w��Fk������k�E�?!��-�l��?���4Fybsrsrbcu�Ȉ70�Z3��]�r�5�������N�Q��\�<���V���ȵc�����۽�+��<��¡�ӦϙY<��F�O�F�[j�Q�.aC����w�����]��0F���l��X˕����������T�2�O ����Z�X�]�8�e�	������S��Y�0o�f�5~���U��ѻ�]�h�'Bi��z���N�N]~�M '�|ҼZZ�Σ��#�Tߡ[�s�(Y�n��7�X����yoB���������-��B��}�%���>V�\����$eki�h�V�s�me2B��ll�@���˅+pÆI�ip(��ϼ�����M7;�:��\�4)U�:xŊ7���Ds�m'^>ꢼo�b�iv|_�F��kE>NQ�4̾JܪܵIjj���Ճ��w�H�50�yom}��ysH慫�hIAK���緘ʂ�@�?��E����w57>��Ыv�E��(J�����%Gf�c_W�v��M�Ɲ��;�j��X�λ%*86�;9~�f1X�#��y�)]U��KnpI�R�|��� }�1�J��9u"�3��L�Ě��jl��$j
�����8�w�����8�G����MV�g'j	���r���&J��'&�h �o�J*jō��PK   }Q�T6�0{ { /   images/c51b28eb-c857-4ce7-b81a-d633a3d7e747.png L@���PNG

   IHDR  �     �PVo    IDATx�	�,I]�U�U��Ww�~Ι��>�̰�* 0��p�EAQ�^��z��}W}>?��wԋ(>D},*��� ���s����]{eVVf���#�������90H�铕���A`<n��ݰ:�t�������꣜�=�3s����VG}~I��ԗ���_����X�K����e������{m�2lA��"��(�B<��rFL���8"A(d����B�"�R>�
	{����b�o��xݍ.t��Y���������2[*�E~���$�))K���ߑ��߷�[7��Q�CFa��&�(�[{�dD�\{��K_Ku��#k���d�d��^�u�ԥ��:B�>�+ʺ��L�R<q��蒆u���7ц4ѥ;R�]��ߑ�t_��G���\�HQi�8~��P�z�{/����ne�^�����S���~�tA�y7�W8Nz�f�У=u�Kt����j���T�%=R&�9��ߑЃs�8��hq��2.|��C�n�?yL���<^�/�׽F������+u��2u�[�v��d%
WA�Ks\W�n	��_!��Z�N����>n���Xle�lu�z ���E��{��jr�"��+쵇.ȻT�v�+*W_�F;$G������(�:��b��vC�'�����l+�ӻ�xb�a;����m�NФ�<�@�ʻT��P8���o���>���0�z�E3�\Ԍ�v����p���g	B��(!5]�q]^�i�M���iEt�����"�G?��F�P0���A�k{���Z>�g���-W����O�9U[_��՚���=��[isշ��7��n���J	��P�,���ns��b1�I �0�u�
5Mb�a���V�"��F"fh�������f5E	b
\�Z-!ON��\Rx���&D�F�Je� C�p*�������}�{����X4����xڊY�*��vHU��~��«��	?0�$5Bi+dm(��ԕxk`��I���Ӫ�_h�:ҬSRlO��M�IZ)^�+m�dsItL�j
|�A�Cㆽh��}�%�1����u��������ז~������a"�58'X��!3��~��'&Ǯ����H��+���W�,��BJ�Ѩ.o���/7/���]�n��x��G���?|�Kw~�q���d2�ڑj��(��f��9�_n	"� {���I 3cd��$�������-��\,b�[��3��z�u &����h�uG�{C�N���O�K#�E�:H'']У ��L��Zl�E[{�I�Zw���������'-0l\��C`*0��:@QG/b��t�v��9	�N]�^��1I� 4=7K9r&j�by����u�P���a��A$yjt��sa�d�r���H�������?qq��6����ly^�n׼�cG �� `�Հ:��P�"��n���FŌD� &E�F�����i3�m��@w�@�n�à� zӧ<��{T������Z��=����>Q0�D�3�[|"i��o����=��F¥tl>����P���hD�h��Rw�A�x���^���c,3��線`L�5Ȗׂ�X�߼���#��k��� �P/�!�4"���:���Ѳ��g|����_����g6� ��Mp*��k~:��g3)�S���Nӫ��57��B2�����x����ut�n�7���fe!�M�tz�o��]��A��xP<䰎�^	��61���P��M���������'� �#����V���L�O��vgkp�JR�<-V<"�0�mb��l����1����f!м�E���6h���F����M��~4��v.o�t�5@@)2�V�@�^.A�h�����w~�G�~��^��M���v��-+X4]�K��8
�"m�hS+���\vă�l{��,X���R���0�i`b"#fG�E�u ��hLx���6G3,�[�v�H����ޭa���Ԧ0T4�)����`�l�c���;���;V�-�xp��r6���7���� ��8kr�LA�lk�#=�i��
C�d��#�09aR��O�L節++++�Z��w�5::r���M��hYV?A�S��������|�����B�0�G>��;� �L:΢dah���"7o�2�|a+���cɈi�맵$�ZJ:���Ax��pgCy�]��ݦ=�a��"юt�O�W�p��'�e�O��!\a�,�ȡp�<��z͵������]s	'g;<^l�}°��ֵ�H")���8N����¹D�mD�_
�X�p,Kg��z���T�V[��o\y��7?}��]��{#����/g%}��[���گ��W�vw�^)6�2�La|�v�T2��N�C�d��������\��'xn��D.�ɏ%YGnd��V����2x���*�08�/}�����#��d��aF����s�R7�j�Ρ���'����wPZ�F��>�ȓ*~���������*�����W�K\"�Vm!�,o՚���p#��L�x $��:��6\^^^]]-����8�w�0���d6W�	(�|&;5Y�֗=ro�.^�k���+7�x���H�٤���钢Yi��9B�9����l��x�\v��-�^.��3�'��ؘ1��,�E�d�rzeuqa�t˨D�Љ�a6��A?�C�j;v�aׂ�s�Lv�����t&�f1j��W��휸�+6(��4Q֡!�_ݬ��+����Rj�xE�Z)˶�H<ƭz�	�Q�i�� $���S���5'��P�����36�$��+��ģ[*�����>G�@���Af%�R��4%��|�h� o"MX�="M^6D�hs�:m�50f���V����#�����ﻦ�}e�>��6Mj�cs>��H�Va�&S�Y�Z�F̑l�ݮNF[n���{�����t�Q��n+7۶���[K��'�g[�x6aeWc�h�����_ر���J����ܳ����y#���v�������T�J%�c���5�ż�A^�;�TP�Ї>q��ii��Z-(��hԛ�T:7C~�Z�?}�a4sik���hjt,7�{j6�����y�UGg�Б���B�'��ȏN�V&�!�a����BvT�Ff�5D���.Q�?��p�p�.bCm&�h�B~�hذ~�0�����# r�Wh��|�]�e���#U� P������@V���2�31��"e����+=e�5��)?�H�B~R=�}�n���P�Ѐ��K�i'q��m/��@�8e��q��u*�'�:$N�ʫ�]q�~�ˏdS)��ٶ�!�N=1K.�} je\/\,�V��MNx�yͫ����ۿo�m����x���2���e�G�BMY�	�4$=~|�c��+_Č% =�P&���@n{�y���*���������7���!7�t=�)[�ɦR����}�|��嫷���rqծUw��K��w<ٌ� �x�n,�����
����' (1H�C�>) ��B6:�R��D)���v���L����*��te�uZ�C1rWޘ�V�TB-�Z���)@}� �e������x�s�����-p�`0�H��y��",y"A<;v��fm��w������׿�U3��z$-�t	-O`�T��J�������?2wf�أ����+��1s�Á�p�O|���������"3� �erQ�:'�e G~�7��؂S"�v}�#��V>����?���&&'�`&���j��i��|.b����w��^��/�ǐ����O%d��e�M̏�jzj�)�?�܏=^�V��X6��H�"�CDDwR�R�)�R^�DA�n2���R���(�l�L3iAf�aH(Ey�����&7�(���4�y=j�����!�#3�:Ga�L@x[&9YqHX��IE�q+I���IR�B�nk4�r�5�D�?X2.���v|����!Ah)9u��ض���d<����9���n��w��������4��t&���d90ڳ���x�E/zn&����G�%�j���B�������4�Lv��� � E���V��]�T�Í �r�X4~�|��� 㹕���,�İ(h'��F}y��c^`��/�����/�r�u�(T�B��rAH���r��!@�h�g�r�����3g�?\�ۙL:�����͒���c%�R��`E����+"�9�)]�6�t�%�9�JY�d�X�@��VE�H�m�������?�L�@/���6��H�`�r�t�>�54F���}LhK��-KZ��R+)�h٪��U���خ�vl�ap	(�k�$��f�V��2��|zuy�����Л������_}ֳ�g�>Xz��+<H� ��fӍǢW_}��W_�R*?rdyn>��
�w_x��GW�Wn��i�Y�i��mtQe��������l�\~
�3��?��'f3����k~Fk"V�,���ܩǀ��������V���r&�H�P{"��2
���?��'X����_=9=��~�?�9~v�|�����"��
�\�'��Mv1����S�M��&"�� >�nԝvPq+zf<�,�9齥��$����h�Q�8b4�s*r��:��� ������4`���,zDV�ދ�>�n���P0���8� `��H�R�=}���[~��~�W߾o�y4l��,��Q��2��V�r	y/������v�׿�/.-�ݷw��@t=֨��q����{��et,�#t[�l<+���W�A:��E_������G��1BV6;i%� qs�,o]�&��l�[�g��?�J��Rej��˕b$J%R��#lа��)0
�{��je�0��>�W~�?��������Ri<���$!�e!��2yv-h��k%�Y����m���&4�axí�_��F��[o��kީ���:i��P�Q������g#�P��b4��D��>"�6�F�`�Щ%���惯�nl�[�{�zd�EV�C�Z��a#�J-��5ȷ���x�k^V��J�2#\Z-�G3����x!�D�`���1��N9�\s�����?
�v�w�\vM"�Md'PO�ҝ_߻o��_�B�����%�q�@�(n�N�������_�vw�E�0�2��4��)b��~ear��?��XL WI�n�z�Dr��\�P�
0�l�1���|n~��������O��/��]^�/L�J������4&?DY���h��V��a����Ukۮ[m������˱S���=���#Ҧ��+j��H�L�NĠ
ȃB�q횈T*�6aZ�_�2�@Q��4k�2�]m�m���XtF�E�\b�"Q�����"a��W���~g�e��l�4�{����bI(2�8t�԰�#��"��{�������q��C�r��+�������c����{��/��禓|�a1���4��+���?��j=<1�/��,�	��ťs�,�A@C�e��^F�z <�	"bp���ZA���� �s�===�a'D~�~�СS���ʞ�T�X,F����IP�:�Q�򼮺Q_T��(T�)�b��8N}e�bE��g��� b��ُ*�<O�b�C��'D'�����	t��d��LDk�]CP�-���r��b ���,�C�x�Ş�/�K��GϚ�1��Z�D�^��ZZ\��۽���w�����j{Z���A%�]��u�vff��++�	�:ƻ������;�E�Y�Ht7@��e�`9O�8�*����}�{��u���]-aB�L�:�4WVε��_��7n}�7�@��%��Z����;�e�Q��V�4�oTʕ��#��׿�'����D�����\��T'�h��ND���D�ZNgR���IZ�x��?��/9U�i6�'hCR⠩���~T� �׬�8y$b4߄v��_��4�������� �~�"+���6]Xb`u25Ѷ�� ]V�DJ�/F�BFi�6z�����~�_o���$b�����r�'X��w��>l��v\D����{qi�m�Qn~�����=S�R��U`?ht�B�^�B� _�uj*�<���ר���A��G4�Ņ��y�G��k������@g3V.�T�ъ	7�V��D>j�I�RįO���{���?��[�5:��+�d��?����ALUu !���jd�����\���#G��
���L,��n������Z����E��n.7��ڳ^1�z)71�]?9!���������D�^ k5b�#�s����W�XDR`�מ���V��;P��R���#�Q�r����ӧ�V���v���$��=��jq�0��L!�hH����/&�T-#'�a��[��-�0 ��]n7�b��c��[��������~d`di��?JN ɣR)R(������l��NE_��������ǖ��kK���m�̙s�S�up����/��d*Ui��
�مw�����k�����=��d�!0��I�\��Rn��ĳ��<V��|�3�����2�^nAW�ڭ���.���GLu�KЙLJ���F�N�޷g�e���������+���M�M�Y�<��X��\�?s�y*nœ`$�-cm!�+�/\m����G�P~��)ױ�����|���>������F�F:m<��7|bfze���KyH]ժ�Dw�S�ۇ��n�-� N��mpU���ܽg��/y�����  ��R7R{����of+H�(۶19}��_{v�g)W��S��X����N�z�?c�4���$D������Z]���1tVKe�DãH{�]�lJY�
$D����V`�EL�iZ�80�o�����#(@}��@K87�N��bC���5�4�N�(.' \�Īa���,ޙ�qߙ�}�{�+�p2�/L��i$-�N]\\4�P
�<ZH��9]�\ȷ��r�,��V�����࣮�X��կ�s��3�Ϻa���^�7�M/�.B(ӀǦ\RW�`;l��v|�-�g	��Y�)��v.�,4�hd 4|������4��EOX��G��0Xs��6��Ͽ�>��3���ꃦ���D�������_GF�VΡ\��0�~(���l5ab؂�5~�0��ھ�DE>�F#J	�D��<J�Y7I�r�sEg���������]S��$��k�E�2ȗ�p����p�=ҍb������m�өĢj4D���['��=}��H��$�u����f�i���I����S+��ü��#L���D&����r�:{�\uu1��y���~��u2�*�v���9���H�D�#
R�%�	��o�r�.�M��0�%~�h�P�O��e��P�5�!$I4Jj��6|6_TtLӌ�r9�g����RX�(�o!�x���-,��C�������Q e�\C@!I���Z�|[��8K���_�kL�e��ѻz��:�z��+9�5EшT���LNl��h��_�V�qh�u�̓f@u����df�� {Q���3	#��z,i�\�=�p��_ͨ˾@�f�v�
6�t��]��>=pK+'�d��1}W��v�uc&?�ctlO25u�}�>���a4T��}���P��d��V:�dne��D�"R)*��" ��.9|�a��[��Z �c������p�Hi��R�"��/ �0R�g���$�F!�'�Z����7f,�����h��Y��Ђ�����֝��L!���	u�3��N;Q�GQF�D�!N+ڨ��JE^�%�� HG`b�tꐾk���.hv�b��z�T5��#�w�Tcx(�;�r(\j|���%���D8�W��n������ફ��Y\^f$Ԛ
c9�K6�:;�
���o����>�j�..�M���^k�	�����v�O\ML����{��ԙ���|�^i՛��Uh�dr�/Q*=/��j�R	;�&����`8�V�ݒn�n��v\l`����X�!��ë7�lRi���P ��Q�&wb�ۉ`0ZQ��-v�d��[C���\(;� y�p^&��2`��*4Ӳf����6��8���F��    IDATx6::��xٞ=+sgw�G���𱳪`a�!O��!RE�D[<J��-+U�S"a+�H#7MXf+ix�����I+������W2Y4]ن>r���)�����T�\w��5	sE�����GB����ڹ��JdR�V����F�jz�b��:����S_OZm�RkBZ��.�.#�f$V�L璓:�����f|��c��T�z�������U�<�g�U�Ӵ���E�;
��ʹi|[hZ
�V��V���#����Թ��۪zVSJ���+^џ���k.�:i;_M_m*>M�Ng꒾�w��ټD��,��%�P��Ň�(�����b�ڒUu}��[�[w�&����9 ���|-ЬV�8�{n��.�I�,.����"�������z��Bp!@��'pR+:2;��Ul8��k2��j��2J�4���i�qǮ>"|f���Oҙ��QH7��Kg�x"'&� *ӹ�Zy�m.X]VJ�Ȉ<h7�b��
VR�!tT(��.stfz,�E�y�Ch���k�"��%��I�h��������! N3��hOà$<I�m\���a�bW9|�:1�G�_��f{������X<?���HQ�8m+V�&�.A��͆h�.JH����Vm�4)<��P�F�
n@��]N�[��~/[{���V*�Q���[
�OtQG��..��.(KV2<־�~��Oc��Tk;��p�,�ڨc�]L&��Y%�ƨZ,��J��S�l6�#3:�P��=U�@�峭��,iqhyZ�F��lm	>�c���j����ۂ?
B^�����4|���ÇW�/�ĉd4�4&)y�T�ۙƹ!��hG�&��Ō�_��m���{���م�5ޥ�V<��N�1�+%���S�Q��HK$�o�k4�-qD��v݁I�Cv��(	�*�N �q٨2��޵ǴB1c	y���e��Vv|tb$�O���NzN��+���-� X����U�#��	����/����ˉ;��G�P:���	u3���]�U)TR�^�q:}7�p�U��!'��V�~�Yj�X9\�o'S��+c~����
��YSѪd�+�t���!w�u6E
w���!e��4��O�KZ ���b�N� ���Ż�z��]�2v��zlt��X��!��\����Y�^苸id�ð��O����9f�P�!~'d�j��<�R�T^"���ղ=59^�ԓ��Ǐ��{����ί�.�K�N[��ZMv�R���J�8��TN����(�yP��Fc0.��A��S�f1K �������Ga	�:�G.$HY���I�F�(u&���7��$LDc�t�<�t&:R��s3;F=���Ԏ�di���}�0�A�(l�֤��6��~�M��g}����@�Y)-3��ڽ�f�
�&�m�`�TD�-u�WW���D7$��\>�ѭ�t�ԧ���A��2�뢎(#�&�8��
%e6�L���k�̈́��y�֗�G�tzϦ���Mq�߾@��T�n��{{%��������]L�Ox�J�o�"j7�^y�{(8�R���=G>���7B3��Hfd5u��G�C�7\��^�P�F:&X	����&��|6ިο���}?���7�
� 4�bdF�`��GU�'��½J*rt�0�G�����!\YΛf���W�NV}?�Y�f\R�g򒱤�䥴�F�n؄��اc��y^��F��� O''�ʭ,..�����D.�t��P�Ie���p6g>t�[G��1�[�̠�:�dvT|Ӻ�2���l�J/����ʭ^���C:���N�ݻrGǮ���J �-���<�	27�Φ~��.�ϲ� �]%�/�	�^]8ۘ޵���{R�n�����Z!Uʵ���O��-�bO�&>hٞ�hWW�}����~�ފth��z"!�`ܢ�}O}���D+P�;5��H����}�C�a��d:�ʲ*�}9��w�5����피W�I�K+��Uʋ��H������?�3oHGs8͵�ڞ2�۞SwR����ҕ��۬n��z./X����z���5��x��	cQ�qXY�_Te�Ee�K����D��j��%��G�=Z/b��ˋދ�F$p��j��������_K&�s��={�\\���Wy��v^s�S���3w|��w?XZ)*�#D{P,�}�_���@_I<��?�(�+�D'eS�Q
���z����vk����/�>�V���jҺ��H{�5T���*b[������P$)���ʧV�6P�.�x;������HO&�&v�-�������^����ޝ�[2jY�	�͇o�+�J�cg�u�t*I��������#)�ht-pJ�y��9���Rl@L��4��ln���S�ڱ�'��W�����x>�ȪQ!�Ej��nO֥��.PJo�	P�Lr�O}��?z�`e"791c����G�0nU4�m.��(���D���kĔi����\��3��v[e�Y5B�J��u�2w3=�E�t��V��Ri�\^(W�q��#�#�p]�kh��#�.OL=|��1������]'�bN�RGO3ڶ=}��B���NQ�[wƄ�&�ꖂQ��[i�u����ڙ��n���MO��y�3����/����\�A��$��������<���RY��	�/��/�NP� WO6]���z��AK���J�:4�b����Tg'醟^��O6�l_~;[��1��M ;�YV��K�`������o��W]w�^6��� 7Lh	k��UP>����0N�a�������:ۏ����0jO�&T��u>�Fu/���!4B�K:.��-Ektl����o�����}������:�|,���T�B���Ĳ���5O�-����S�O��<Xo4�Og��tVzo��=thF+c�F��p:B�c�ݮ���`��0�8����+�x
˝���z#��_#�����D�1���WV�W1rB�8���]���{�[qi��1���$=A)�P���w����d4��dߩ�{�z���|W1h�s(�����sdӤ�������x�Gi��l��68>�������؉c'��,��,T*-#�����>���+�G����DcA��w�'H�B<v|���_:����'r��e�ؐ�kd��]?��-9��PO�C�63��QV�ۮW#fRx�a�w +˳o�?�+���g^]%�M�uY�s��Qtr��������?�����0A���,�ʬ�VQ呢�q�#]:B�7 @?
?L�@M"�����ryrj��N�;�ODC�8�4�F���x�����c#��&rll̲�!���^-,�T�}|�|pL<���;�y�M��'�Iӊ��H:�YXX�����{�����H�2��dM`�kZ�#���{"`C�����P�"z ���Ά���I��<ZP����^���1<��E�H4 �K$�GZ���x�hD#%�s�@���2�AJ�����ty0��$�|Q:]�F�@���c%Q�ل>�I�4�!'��:�l8�GNh)�
t]y���h�%߄$��V�,L^��3�r�y�3�l�L��3���zG�����������a��|��l����ቪ&�%v��]Z^E}|l|����(.�{��͖_|�ς-������a�\P:��.R=M��q���/���V&R�-�N �����n��fj�IR�D�����.������@�(��M������f�����?�������_�֟zL{$Ꙟ.��7�����oz�;����!���cөd�Rs���2��R=^����v�tc~xC8���H���_�:�ˍ����fvL��?x����P�Qs!{��? Z�y$�j/���$~U� �M�e�pD�����;?�z���]�������	 �#���6D�#��H� 8>)%��;(0��nh?�Fs��\���@���ߔ�~�A����e%��g��<����hA�O��������ݠl�s�r�r)�a�lD��b��ve�qY:�,@����Jo������£��>��>��,F���O�\cՋm&�IdF�iL��� \*�FM��DE���<�����>���+Ҥ��QQ��J�GŮ��i���W��o���~�U�~�����岗�占��4;�*0Ξ/�����;�<|�d4>bFS�zk&�sB�1�/�����T�h�0��r���2���k����y0���ڽ���od�t*�
	#r|���C�։�g��o���?��\��Fq#?�뜃���4x$@���q9%���^-�����4�m��O���[_�"+��aŚF�����J�} ��{�#��� PL�^�;0�JtC#H;P=^C��͌ǘ�k���ZĚ8}��
p`�*X��Q�����)��
 �1ϱ�9,��|��S�@��f%[ۑ�`�S�Y;��E�I@�{Є�M� y�I��"-�]BZ����Щ���8���=
�PqEx�<D��l.e���N�YYD^`%�/�����E�.t+�=<|/�Mf�pIE�KU�4���u`�lEc��y���!��+��n�Ü�d�U�2��T�4����zܦ�I.�H�]t���z����RzK T,��{������|��C�˥|~�կz%�@++2te��t.�Y�{�o�߿��O޾���7��O����"��%�|P:j�x\�zDq.c]��f��3Q������動)�%��_��o�=YȃSn˙�upyyYm>�TʱJ���ܢ�MF��t��͖��P�JK64R�x�����o߾bq5	\���Ď���w���o�{^h.�tB�x^"�d��k�y�E��R�,e�P_��ƟnDUV2�w�(�@(��m9���'P��$0�BA���H"/>�By�$���ʫ�|#� ���z���t�8`�RR%��P'�a~@�	7W�&������^.�jG&\Q��V�kc7*|�8�� �����گȝ���*ԉK�Z>���٧C,�<\#���:D�`X��5�)�<G}�Q�*j�V5K���,�D�G�@��$q�Z4Ȥsl��\����ذwp���vJOb]!ʳ����C�~�oP=�t���A$`���i���vt���/����w���B�)!(��P{͠�`n�?�P43���F�`"
/3��ҥu]���Ou-�wc\nh).	劄��t^$H�F���qF�ie�9ñk��-ҹQ�\���!�pE� @�ʨ���b�L<�e���FV��qc��Js1'368��A�gee���HÁ�ٱ|l�����8|
�q�2���#Vj.��ԛ`^6T.jT�3�S!��:O���=�e<k��V��<N������d$�`���oPHL$`|i�aT��i�P�7� �����m*��ix���o�Ԥ�	b"{��b��]��ײ�mX�H�s$����A/�μQ�&���<��i��er�����AKV�x4`E=�<��K�U�1�q)Ky�5�Y�`Ϯ��Sa�"4mKŕ\4CeU��q&1jV��5�z
] ���
	�&ցTSu��'f�f��Z^^��
�e
̦�Ґj= ���I�(�S�Y�O��- :.�I��C],���Ǔ�z�}v�je5_\�?f	�BF$�*L6�����A�'F6�E���H�_�Z�!����Q:n�'+N�o�e�ߥ��c��T��R�.5rY�	�	m)|�P;��
�IdG�c�)�e��%������N��m�ľ��f⹄��[k^�D�0|� 1�x���J�@2d���R(�b����t*���Й�� ��'�VHW8�H�*u$��C�Fԃ�8h�gQ�(� �L�k6f�Vc�|:f6^Z�Y��-�Z�uiv��]*�GV�-_��Js�sg�=�A��������W�r*�-�g��Y��cq����)�(�&��G>\Ă��d�"k���"��'�|p����`����QU*t*]�Hvr6�Y��C5h72d
��l� v��7��g���?��>�J)�H���Ru���H&18C����爁�U,�p�������v��n�����r�Ѧ���&�X��_K�7V}f-�Ҝ�Ati��^̕�C�2�3|�{�⁂m;K0:� ݾD49��&�2ɧ�	���z#Q�b�'g{k���M��ئ�Q�2�����7��Q����s

���޻��������C�,>&͙�8d_�ZKg�-f;5׵�����q���rP�c�Ċ�ݔ�1����	�����:�C��"q)8j6�b�T��mgң� ��$xX�#y�D"^B�@-����	Յ��S@���U�$�T�K��V���X�.�_����Y����\�	`A���1/p,T��=dY*>����˲�C$B2c%������xnC���s�u��>+k�`�0_F�t�q�Y�%c�Eg�$���I>�f�PpVk��H��*&Ƭ8C��FF-�x�Ċ�dJ�Q�."��Fx���DEc|f����?���?��0$���d��**O}��hO7ċ�]�u�bО�"��wi�N&�����|���������"L�����ܝ���Q��{om5����3�����հ����Dv����	�����it�`��M�'�`�����1�;-�����fa��t�@�uC8{����$�M�D-2���_*`#IA���c�U���R����uj}�`�*b�IGFc&I2l�P"Pl���A(<�T�\e�0���b���B�*ῇ8(22�����v��������"?�)���j)a��+�m9iح��<�P"GEDE�FC��-[� B� |!�����>�J�R-5)*��8��\�Y��$`��x�����9W��91�+�F<�"�(�[��\9ضDQl����K_�b�_�g�2�W-��#������Z ���Nː�<�fX;C�^�k{�LL��!kO�m� E�	O%�&}@����o8���)����=��|j�U�ך�痗��Zu`yxPz��R�F��)��fc�~�-cc
���}����_�����ܹ#b��� Ȓ��@�s������p�%M����y�s���7^w��JE<[G�I���̙�(�Lc�b-��V��]J|-��r�G����oN���<�
FP��%T"�DzS,�����b��:��t��2ng1�k2����8�T�`rf=vnA*c/p
C�t��c|�ʪG�]�?�^ S��.{#�N�f-��6!Qd��a��t�BvJ5�D�VZ�'�1�:,��F�A�X���|�Ʋ�������:t��ա8Mv�N�"˜� L���MѠ�ny�u�Pj�n�j�f���H#�(VVµ��8x)#��qۆ�邉�xC�������Y���8[o�9�	��-��P�R�г�B�D}T��X��j��IJhs\�!�e���B�o7�����7c3r��3�B�_�;KK�z����o��G��|	/72������=���Ţ�̎R���(�uU��	{Щ6�Z+�6��|��{��W�n:5�f҄_������?�;vJgi��SV��eY��3�� L��][-�!�����ɷ�qz��^�Vu2�]JN~�w������J���1ڢy�6J<j5D.8E�	�.�ܔNe��ji|lW>ϲ����ٳſ��O�ȏ��0�:[;����3]Q�%I���r��(�.&����2�A,/�c6�����O9�������č�_��#�Y��� \�z�����Y	���׋W,M)�|���Dtg�i!��ר���`�`��t�\ƈ|�V=]I/k��B�+.��)ဠ+8��a�a�C�X��wgߥ�6�$��L��Q�_q��zL�N
#���W��N_ɝ{�-�l�c�d��:jw�=?|'�[1��z�P�����-�_��R�Q�9������A����:��b����9��t
$�J�%x}��=��-���@T���l�#e�n�j���JE�cW��ރ�u�..5���3E�.x�%�-D.�J�����-������=ik@��5��h���V5N��fܟ�؈T    IDAT�aJ 9�PY�t "@ݿ�v���~�N�m��Pk��P��Y��x5���Գ��l��S�cfd��^��[�u��׿q̊����xH��9J�8|}�t�(�Y&/aB�탻��Ν;�D��\>�Œ���ȁ�ҙ���*S"t)�p�d��I��"Y�
�Z���;.��� ��F�vuY<Z������� K��'e��s���y�0�YȮ`���ϋ�ٙJ�gϟA�`jr'����>"���:���Ba(��X���y;�����x��%��:���8 ��2�:#�s���V�|�)��((0��mп���m�Ű�/��k�&rT���JCl@�z��.�l.���Z����RM$A�%��G���_(r�b�B��ݧ'��;���W�>�����{54ۡi��2�¾�k�q����!�K�u*v��Ë"��	�ڐa׬��hi�۰�QR�,"�v!���I�)#�f�����9$H�OD�φQ�}_,l7VR:�z��F&�Pl(mFA4��  ��x�>�Ж+�4"����8�HLyJx-��>!IЂ`�R�hF�[�Yltj��je�kű{G�\�^+��V�[���pš� �e�	
#�T�oԗip��h|cuuE} �քU��%�o��&�5&n��B�A�B˦3c�b??0<�$GP|B=ү9j�eeBY�\�+:(ɤ���(܃�a��~vtW6?���*��F:U�XL��D�����W}�w����PL�)��I����� :����U��˴.��l�|�m
#HtsU����b��J���'�Q��/�^_RRy����?����]�G���ݺ��P|)i�G5'��P�^ҫd����6;l���@'ȳ�˘�G�5G�~��%���:{��k7�q�L"��y�u��s-�ϑ��EV��Y�����H�5������3-��ݖ��W_R�z	�%���}E1OQN��k��y���u�Π7��Q(HC�PC�.U+�Z��v�͈[��Os)�H%��'A,�X���y�e�0t���ܞ��^<^,-�q��eS�R�R\M%Ŋn[2�G�M��<Α��<؝�,$?�C��x

�(�W`F��z�_:a�p�Jcթ:݆��<���g2�-kF����+R��p޴�+�믹��/x�W�b,a<@>,�͠k7U�t�p��W�����P�8nY<{�������]Z*2��2A���TZ��m-��<���^|��u��8`��_����|	� N�(#C8˗''iV���BUaî��
��|�o󑯧:����QO��,Z��t���2�X����V�L_�t5�:-���wTh�?�EY׈,Fa�-p���HV����L)���o�����f��_ݱ�=5Q��l�g���Y��1gj�J�!�!���V�����IA7�꣯2��rYD���ݗ���Q|<�LM�Z7�-�F��0Ƥ_�߶�֨�M^��{�W�hR�=�E���� t�<�/�;��,E�x���B���c�p�װ1sb���['ru1 3�|
��h<� I_^-=��Cш�ǏG��q��E����)+gFj���e�$Y`A�z��P�WG0��2l�q���-/��J����4>=62z����Uh��tŸ ���\$U_ݶ�'܄͊�)xB�jb(�g�}J�-��_�����?��O�Mk-��t�������zKШ-#��'<�S#�d�Idaٻ��>����<en$�ŬH:���D�w��BK���Z�C��EV9b���3q�_6�bzk��2;�0���	���L'���-�l<jbs��%F��jD(��rBCo���
� ְ;�����J�2p�Z�Ϣ3��E����2�	o����%�J�uM}�q�X�g�v͉�������:�wW6�K%F�e!eZM��!+|E;�<+k0�œ���ODC͉���L���?� zA���;�%H$�R"0��T��1�l�5P��W�n�~7�~�|Eq����"q.�2ƥ3#(-,���wd2�����z���G'#y��*I��S��N|;�x.r3e���8�Tp���Ӌ�Gq�1;��%1�����#gu?fAԃ�b4�M�BNED�v8mU�� z�СCG���iqanqqaǞ���·Zfl��
�4.��O#����\��I_���y��Eဣ����! :�{Lf�j�\^e�(�	U{���ࠚ'�#"���X�l��~���ТE�7a�b�
.�ج�	������c�Z+瘇:am֔jwc7��j���;ks�]������/�1
�!+k��ե9�LO-Vti�X/��n-��ƭ��o-��x6�冕�A��t�qX<��!��!���[�3՜㲳���a6���ٽk��3g��]=Mvf5j:�R�?̿	.���n���Պ��s~2���z��n-0S*���i���Q���ʱ�G�L�ɨ��.i	�-��ͷ�}�-��É�����[.��'����Ę��<�|؇ߔ�""BS	8��d��j"��&�q_�4�tG`;Iaߊ�4�]V�L�}�b��a�D[Z��9ɀ1���D� Lr@�ŒЊZA����{ф��E�H�F� ��M�z�dC��dEL$%�(� +�b�C�i�coQ����h�H� ��
[��Y�E\� ���;�6�Б(D8��:l;�?&f$FbьkN�M����PS�e�oc+���ͺfm�u�g�eX����F��s���`�&�e�9��C�Q���tX#�c�a*��)����F��t�)QZ�T��`X�� C�:����^-�U(	)��"E��w�\Ħrk+��N�t�zGڶwN�����̣z���%l:Ryv�Q֗�⃭�e&{q!5Ĩ!�NO�=p���~����vO.����Kh�f��:몃{�s�M`e�=r�/��� !�=X�@�d�-�����E+�L��Hܱ=��V��P���=r�Ql��m?u�Kn����1X �fs@G$��_����hX��J��v�\t ��(�(a��7X�������#X2�A+\�7}L31�^��)w>�@ּ,�r��g��^Bs�-j���I.���Y�x�4Z��B>X��Y���}��6a���|�!�k �/d�j�J>7�b��3f�Yff��p�K�>X	K���d�շ
��O�%�#a�k%d��F�	[ v۲�i�(r��,���K�d��+�3���1�Pv��x�Zx�R	�\+2XgTl�4.;e�� 䜊�Hg$s"i��4��i�+��j
���K_��?��[��j?&!��j��1��"�r�L�x��E�&�
�``��Ot��By|�Gc`<��oþ�����g�G�+̚�wX+�Q��&@X8M�k_�����=w?0=݃K�L�tQ��^�9����##D��pZ!�P����k��;�����?�Wx�݈��w���eK�@n���b�^�Դi��,R0jB�n��!�}��o��3n��֗������ӓg�"ڨ����&�N-���3e�*�ݙ>�6�\D{O�8�lD�~z�������3�3���r��ڹ�+�?=5)SoT�-{�0����=��Y�S�Ѭ-���P����"
2I��a�ԯ�z~��\o���H�ٲJ��y��i	K7�Ȣ	9�h��d�1+��M?�h��7�\a�-VW�c����.ߛm����a�c� ^�L�>J"��A�aW$�H#5�;.̝n������S\h��|��1ۮ"�v���y�� \����G;`�c��-���q�N�bc�;����-lp񝇡3�0pTW���Ȅ�E�U~ !�D��^tV��a`�梬�?��8�p��{�\��gްs[�f�֘�ʺ'��I�W/���\���ݣ��.�wWx�})�m���߅�Q�/�˲�̜����E�jĳ���ml�'�zH9{m��N�����5�v���r����Ęn5i#����
ĔT��pa����x��e�g��I�RA�����ǽE
����s'�4OY���6�f�^:{��c�3ӵ��˧��T�]j��<��0�dh	٥�sb� a�􈻡�{�o�[�P =qpQ�d��r_+�a֎dsW^sm.��2����ٜ��Լ�^�0t,#j{%�*�J���-G܇q66��8�!�g��+�8���J�N�L6��=��w�U�Á��`�όF��,"7E]!�������\�sB4��_�S;�8���=/rmܦH�B�PF?4�^��.z�M:�eV4ia>�"��)X�s���Cٶ���t�4���]��@�o�C��dD�K��7I;�{��!�.��b�]�R���7
��6<��H4��A�RzD7H�|i��t�r�*nJ�*�+�d�ݚI'vLό��2�z�ٹ����}�}G߅���]�3	w%�w����qth�C��g�a�Ӥ2=��%�����Hu݁w���u�s-O�$�v�=k�����6[oe8{�X��3m�hjF8s1�����1����e��qm_=6I�!�'��X��9`��f��#���2�a�h^t��+�1��O�4�b�$<z��t�#���]�&�r�Đ��pP�#��C�I�9��^���6=�Δ�U�a�T,1��H�v���hS��6�C�
�B&�R&�|���^�����l��_G<F��K+���*<w��m��A]dd**EKH�K$�N	���5M�ً�$�{5V�W6"��`���"��#�W"�\jff�t<j�R��CA*�ʺ?:2��mQ�1PxФV���峆"�ZR]�L4�Q�ܱ��sԤ���LN���)��y�� �(���Q�t�dh�ӏyk+
��ۙD~����Je�:Mf���d2q+��g@���:Ω��=���
"P#�������h�Sf�����G���6��"�?7����ȶ� <�&3�@�=ۆ��=��g"�gˤVҊA����<i(t/C9`bxI�+���������'�A�b%w��'e��X6E�l�M��q�];r�.�ѵ�"W�ED�#�1'�":���E����؏J����'��P�x�r]��c��|�A5i:	��Mf�\&�T0i%0���4M'_��\���5���;��o.�xA��r����i8�zU6�Ff	��T�2%�<�y)��#�qѲ`�Jh��잙9�h �������AK��p]�3�a;�!�=�p�gK�*a�	�J���^�uV�8�qg�s����+X�$-L�Ë��?|⁇N,1���,�-W�$����e�;����T��_ ��}�n�og�AE-��T]�J�i隖�_�5�r��GІ�{X(��%Yq��B�/h��)]�A�Ƨ��0E�����
��L,�vha�
Y�&9��FFr�'[��Z,��b��t�
X�H�� ����/Pg(��DpQF�N<4�rz|��STd,`�@镐x��Ag�L���3ܧ�/&9���H���������L˫%�V(@�ӈ��1f7e�a��*&�����W���,V3�N ��Nc"�@s����(z��!�0�t����1��J���W�T]Rr,FVvA"ZZ8q�t"qd¹�k/�b�tш���'N�=s���s8��%-��-ǩ�Q�� \�M���2��Rڵ�Kr6.�|�B7:D�a�Bz]2���ݔj�Z�pW:X��L�O�K��s�~�ޕ�!V������K�x33��m���}����W�փ��֙�ŢY��h^<��Xd���F2vde�A�zX��T]������KQ�71�iX� ���3�|!m$̖_M���Hxy��s:�y��_���J'��2z���s��;>�w�>�|����Jqb��0�SG�)b��*@*.����#�V�]�[��qΜ��Ue�R�nʘcm	�+�b@+��ƞ����]E�GvO���J�B+��)������@�̋���EjK�����a*��k�݀��p6�?0��� `-ڙ(uB체	��n�X+�@�[��px�2�I�CX䗱�*�m|+���H�:m�	� %�r"\�D��@�ؼ�Wa�����h�֠$񄕃%�T��e�6+�&"-� �	�[��a�lˉ�S�o�B�4�G;MyD ?6��_���I���#�?H�tk�nt/��H���Ȯ�[�y����Y�����[�u�5�\��J%�`��<����*�G�<F˷�Y&�d275�{�Ƞ*�
3$�,����t�K�,��_*�Y�|Tv6�9��.@�(G�4���܎�*�
�@'��!���{ <��(D��)����n�:)��3!$~�)^4:���"����L�2H�����\blvA���T�0�bke���J�dZ X�7�:�\���[cC䥀KAb�? (�υ8NA�������t:i?����S?���?#�O�����¹�g��Sn��9Ͻy���x�K_�k��{N�+-gQmA-qk��
�B����*.Jm�����OX7�Y�?���&�Z>a�L���=R��`��:�+�a}ZZ]q[�u"f�q+�p1�k'R�R��0�@�v����
U­�*�򽆽R\Y�L�mۜ�]`M�)$����yИv�{T:�ǃ6��Qo�vs�$��AQ=�+{�	�=s&�ȡ�+���i<*��=��*f"d��d6Q
�8����숹y��i(�|�i���ONӿCM�l��]�Hnd,�H�Ė��*m/��k
�5����!@�	�L�(K�\�&��D�	��0� .5����?�a�{�`
Y;8\n,�*�p,�-&�,&������;q���S&�g���_�bc'[��J�2���L��Lalda~ieuI��XQ�v���zKM��GY��O�o;�7�z�;:�ų*�py�����E�ҵZ6IfN�|k RS��S��ѤG\L�տAp�|�������|Ϟ܍7�899�ģ��#�b7��FB��,�^�eD�P���W,����z)p��T���jBxkdֆ��_�o�JKf|��I�Hqد��f�6����x˛^�co~�Z<y�W9���p��1:e����g���������_�[8��B� ;�G�B(.ڛ�E�Ht[�x�ź@z���t'��f��6r�-�*�$1I�$���8;��`�o�����������O�R]J~������Yt��D��+f�P��#�ǚ*��Qm�����W���dg�kNu�x�Ro���v\6Y-�8��J�B��D���)��f�V*J'�-���߸�v+6)���j����=z���{'dk�Vy��[זY���u����#�<#���F�Z?����r�䣷���Ǐ�񳳳v��5�tʣu�2)j�Dq�wp�"��H>a/@���}ey���-y,�=;���	ї���f��0L2�XCeU�E���`&��痊+'[^1k�oz��ㅝǎ~�K_�z���õW^;�ߑ��w�طk�3���-���F���?8�c'���塥��\�Z6,7�0߆�U�\w,�koP<H���,+��� GNX)�5�9�48�F���Y��@�F0N�����dCG�?2˪L���av���;f�\}�S��D���I�,D�NB���i+��؍����OO�^	U����Eݗ�a�IJU@���/{�<������}��nR
`�EQ��X��_�^�s���W��_�z��#���H�n�RO��i/���k��������\���S7�㿼��l����k��9���0���
(X�:�P���G�Y�W�KtO���S�!�e��p����Tt�9c����{ �u����:��ȁ$���LQ��if��<���c�g�ښ���r�k�ٙ��vg<;�v��%{5��,Q�ER�b @�����u��9�������]���8l^�w�'��?���f��cG�G?��̒H\�'�����Ke�=���VW8�;��re�@x ��R���߷d.���O=�̯����R2��p˾��½�9r����݈Hʒ��Y1=�EՐ��Φ����SO=�7�'��>m�    IDATs���]ݑ�9b]�~�D��R*�!I�Q�~.�
��Ji�*�+�`rr�СC�Ģ}�ji�ԫ2�-$_y��cG�����P)������l5"QT4<����
M����5���1���+���_n�<��XRn��������U�]j��������j�+�R�db^����Y^ZJ�r��R:�*�	�@�	r(�G�n���B"��/
�	Q��%
�e��4cD�U��f�E�ڜ�M��峞T���aN8�	�A�7`o��-}��`F��E>�yU���E)�u85�9I�1j��ĩ��^��@{���0�Jh��o(�Ju����zb�@L�1�أ�$?��P�e�������!�JX?��ݣ5�P�!^rjvf4Y�TSaOӱ�\�#��>��?�������3G&�����C��;2X)@g�
���>�ē������?�D����7����?Ǵ�2l�t&H<��|\D@p����T�¦Pm�� \�;��:���R���ٸ�`�XW	����������-�݅����L<~��xR �=;�n��`�
I��<d�͢)[uT�.�� 4�;Jǁ���\"G]�,�HX�z)���d�eۮc.eq���������s� @�*IN��=C���k�Za1�4_K��Pl���LA�Y�JZ�I���l=���ł�ه}uqg� ���0#�gU�=��~p:ZB�׹��>�Q�D�����=ǉ���d�>"�OA�ß�b��.�Q�p���m�����%���Kc~w��n8�4�;}�AV+eL�|�,���h[V�يB��`�K�*BK\���2������p�.� R��آ��b=��xw�X���Y_*#�H�D�@�H�S#Us뇀��P��r�Bm�38�W��[,�T��`F��8@��Lɳ�[	��"_鲎�`4VrU�!���������$��ځ�&`_�a�k:����%��d�|*a��X�uؠ���rE�a���	�G�V��@�l ���E����lj����][9<-�΢(�e󾑭;<>�CEUq�r�o�[1ffC�+������%��R6�p�,DUV����F:��e2�X�P����@*yph(������p�J����?u6��B�J ���!�8O�5*5�Y!E�J�"r�b�J�i�8Ml-��p�^&�6'A뺩�zm@���P�P( ܆jߦ�ؗ�� mK��􍲅q��}����T/����v�`�	W�^M�f�+ Zނ�k(n��A?���y�e��=��ø�C�	��� `����c��Lg0v��`L3��j�RR�ʀ1�>d`YIB�oB��~��>��i�&ؑtt�� 9�g�Ll 
ہbƓ�F�F6�b��S�xqm�C_��ؘG� ӆ���tY� }$N�g����?��jf#���0iB���u��eƟ��s�"�Y��|8��f�.�W�U浟_:e�%*w�{ V������]�l-ǧ�K�@0v`���wT�~�\>a��J���D\�K'O=�.�>�o��������=����F@,�_�o�~ˠ��б�%U�f�nx!���f�J�p�=
$���"�Ҫ�z�%��꡵#R��o5�J:(	o�/�it	�!�A�r� �����[��^�����\�����?�4 �E*A/F�~��8�E��6������{1���M��!}�pJ�]���G_�3�"~oe5��#�����8�a�0��?;9;g��q�G;!�aeBZ�d�J��C�:��Jd;J1�����������c~f�!���X,�}���2/t�-�'���� P�Z�`w	�5�A#MO⚗�\��2j�`�0 �L�
�ȉ��&���k�A9��<udm��L�V�-u�F��"<�ޖB�dc���2�t��@���ʨ<U���H����:���>f���2r��ȭF�?�XWP��]�`϶}�ۏ�&�H����m��h�l����������O:5��$�(�PS���`��j�S�[4�#N6����q">�  �\IDO�	=����·f!�.!q��,�?����t/���x�"�y�Ғ2)A8�\A���_��Ͽ��y�.έv!5�#�U���p]!M��j���DN���`$���8�ˉ�C��ka�ػ���t"��څUs�Ϸ�,q7=~l���^*e��i��Qw$S�����)�ɩ��Bhp���(�5�ff������w"3���r"��׾���9r��5�y��H��*�%�8!�C�F\];�f���M3��l#SP-��@Ao̢Ҁ~�ӹs�N4q�����$��Y����������Du"��.��m۶)^��:�y��j�(� ��o6�m=;�.aF���0"�/R������q�k}`V�i�Jky�P� �w�B~|� f=%W����qYKLϥ�r�ص��+��v2m.܄#�-���� �j�xt��DghtS C�E�h@!�K։���DƽU�-V0.U�R�NO�铟 �ƿ�(��ҥ��!�aGI|�M�;�hx�V�}�~���~��ڵs���y��`W@��)�.�|ʡd�<��d'!"HSA
�����.�]'Gu��r0��� X�����v���Fi���1w�q�Wf5'bz�p \/G�&d��&pv�l�/�V�#�0�NBf%���`xd�����ٙ�	�'�x��ӭ��H2���Iwt:�8���d�V�D��U=}���O�C�����0F�b�9����z�!�K�*�@���[����5ș��L��t ���S���[�Y�vؙx��fo��`���	Ni�ơ�AV4gm?�yt	[J	�Ȑ��) �#��5�.��&Ϗ%r�]���T-	n�X.H�#O=����L����H�wԹa�!��
m��1X,���22�Opͯ[ť��,Q�N�rY+�k��U���ID�`���KOW� L2�<��H��A�PO�Mx�*�"�"��6�9�#XN�TW ���z��r��Ȁ�j.?l��D|�ԱS����@���WfY��;E��_W���JP���*T�~�݂=5��я�HGf�&zG�)E.�c�g ��wy�0=���(���'�QEt.�ms(�BǪ#�O_dA�7	�?aRj�h7�G�O�"���]��>�����FpGr>�XJ/��;N��>�ϟ?ϓE��%�UW�!�7�4��ȥߚٮXD�@F�L�bH?�add��������!�T����:.C�?�W'�$��ԯH�9�S5��`�A֌0yh���sm�[�q�.ծ3����O�<����-f��	��<)b����<y.�\��F�8���'N<6�)����W�
�,!]8~���cOF�Eo���M,�g�0J�;�v7&���%k0$n���Y�B620gr��:�5J|e��%��47F��������!�H���@�t��+�-��Gj���P�6��!��H�5�ԭ�A��z��J�9�8A#2/΅8Y�1����]��z6Ł[�>h_#��YA����������$2S�d��P��!�-J3x�_�6�z���2`i��/�Y��
�K������_Z�t�#������v{��EX@���A���@e��8N<�劳��kǎ�[v�M+���X1��	v}���Y$��繑 �CAy�(cu=���{V��>�.��sώ;��8]�#�`S�+BW��4��O��:B
_�ͷf
E1��F~]q�ym�+F��j�+<+�o5t]
/R��K
0'f��NO�X����\~t�ޞ������_�i��֭�[62��b�i/���/ν��޹��{?07[���{��G0������YEC���{��QGA=m s��	Ę��[1<5��h��n2)2�����A�DHv	n���X��Y�%B��C��Dv,����*�2帪�<i�IO���d#�����$�{�̾��922Z�r��}d�8�E~�"�H�}�zQ��=Ȩ"lFa�Z־���rJF��47p�'tj�㉱338�������L^G�S�D��������΅9�\����������#c�q�^2R�����;����l�)\�A�����
��ؙ� �Y̤P?U�-t�E�%?i��enV��g���t���j �f��}�o�@B�W���X]���L��х�Ot6�4u�M]��["��J:qC6]`�ѐ2��+��e+~�a����a���-�1�t�=�b�p�0�p�K9��6�A��I&���������;|��m��W�Z���}o$<v�й�W�����-;��������ɩY�Y�0w�XsBX�ꖍK:cG���|��hHt��r��qk,�[�U\ZE!<	���%��#��d�WL���tªzɩ�q!I�Pg�	�Ҥ"5�?�,y�n�)���a��i֢��'�� ����!����Q GG���/\�#��(����Sh(uE��]��G���_�]���T9BoN7P���B��_=���oЮЛ5���F�2-&p�b�3��c4����~�?|�ۏB]@@4�E�A�O6tiP�VE�h�Ju��[�͒�A�7��]�/QO��,������ٳ˽!Z$A�[�2� J~���B"�h1�	(�K	�Tڬ�?���f5/��W�aBuk`���x�#��گ"��+����Ѡ�Z�C���|�B:):η�Y�=�+CD��R`����[����)AfB	��r�t�|H �J!'A�6��pG-$�O��֝.�){#�~t��,���-��⏳��|RTo��'�����g;v��y��ݷ�7[B�L88�c{$��1�pl��??����C��v?vи��h�s�?�ߛ�j��WI��<��)�����������}��[4��3�H5�"��t5�̡���R�`�.��O��q64�؆ȥ��!��R)P>8���~���f�C :X]h�LD!O��BوF�08�q�Hf�eun~�Na ���o�;1>>y~r*��bySKT/?���y�1Y���aµA���!T{9��C��\7�wt�閽_LB*�� Mƍ�0�F�lp9�W<B������)�)��P�R"��"B]zhؓ��O���W�-����U���Uvvo@�G9��,=���R��864�����C�o߿e��s���K�=;��{ێ���^���z�?��'{r�RpA�:���/��;�.�����}ԥ��`�2�����39gN����w���	3׿��I,�oݱ��!��2�Ů�CT=��K/)Ap���������V�!B؍M������z��Cf"l��=�ra��I�� XP&��I�	+ec��ғ'W�xL��*�T-�6+u�|6����P�ӟ�@8���c�����X���$����Lg��w�%t�O��@�^�|"�p=��"z��$��$O}�����ܾ};��8���Ȉ)0qNX��$?��!�9<�Ꝇ���d�:�F��%f�+�<���L����=қ
+Xv�6����<�87����ܽ�lǐ��[��<�T=�⡗�����ȏ����H��\HN`3WN��-���з,��j��щW��v�Ū��h(;���ɭIq`�VLA���Ǐ��ٟ��_=���=�o�9��9H�������,<��� �E"�f <��檤�AL������ݽ=�4,.�/'g"Q��>��?��-#=�b�R�"d���ؐB��l܊r�W���j�A����H�ܐ~B�B')�Y��Eo_�B]ݡ`���Oq��1J�p�^�ĩT�B��:�RF�D���ּ�v��Z����#  lE��@7I��e�NL��Ux��I���_3>|�P0Vd 4�l�WWB��@if�'NfHT���ϰ�� ޼�C�yt�;P
+OhK���S䑫%�Ϗ�깩��qt��\w����0���Scc�#��N�<?7�)W=�����3��D-{qAؚ/w���ڭQ����*��4PgWuX<�@]�	6��C5�������S���Ы��ՒG�=s�8���w�aV���@��(�㲉
�p����_��f�{����x��Ƹ�΢�SIa}����F6o�2�!lt��=;qא��X�B|��Ti<����F��9��=���)�(̨
sU����d|~~qa��\�$�
g��~"TA�Y����T+�8)�ނ�>�'a�U���W�t�Gݠw�	�l� ݧ� J,���}����'hL(�� �C5�d���Lʡ԰�NC�q��Z�a''���8v]�ˣb{�)0+6z|}C8+c�0Q�]�>:�1\��s�=�X�WD�"�����A�x\>�pW+y�����c��1vM�j_�}?R��/�%e�I&�V�(��Ysڜ��s��^x/�Z�oSgdX�JrR�<�}� �~��T��D-q,�� ������~;66�]�x���	�0C�	%�g�J|!�bA�;��*����/)D��V!'{9������]�b��,bD��D����`���[vHDX��"!�eV�Fy͈�Ćju˃:�3�� 6�	��aW��&Ew=p%?Qjںu+�mbb⩧�:�<h�̙3SSSd 3#F��f�'e7M9��"���M��w�/6(XX7ͼ�3z�"�G�NQ�A@�fl�� gs$>��`�Ή�lG��V��ٓ�X�rG����W�N𒚷׼5Ln�¶zeI,:wjh� �	�Tm�c��B�V;��v���5 Z8�r͂[G�L���ž��Mw��B���8���0���d|���?�����a�/��x:�>�K�Ǣ�σ�7�W5�t��x ؃�ۯ�:���o����b	�5�X���g����J	��J6���:�$"���F�`L"̩~4��Xt}�*�J�'*�I���e�"��X��sc�/�v9B��Y�zgFH�'qf�$2)z%����eO~�X��u�N��h�HD݄����k\v�+����i�N���ڌ2z�x�<|B:�D�]O~�޽yO�0�|��ɕ�w]*0�� �*�6�6�f�Y<�[�$�U��U�N����Q��0��u���kB�ßJ����@Ѕ��	l ��l�qM{�qG N"� [�����d,ڇ@mۻ��[�8y|&���n�{�3�S�P�\�ypF"v0�r��j�V��#�%*���[�p���] ��#zC�@8�_ʥS;v�ڌarܜ��L�$St�%��bV6ą�8 l��.`	~%Ǝ4L�ő��$.(��3	��܊(�se�j��W2)TiR@j�h G���H'�O.n�u���Anٲ�%8�-��'\�[�(�',�g�y�����9#(;�:�F	�k��j���'H��|J&&8�Қ˿b�Σ�Jۅ^�+��y��w#�Zw�q߼4�s=~zbށ.Pئ|۫Ƣ;�D����6u�墭��+��/'�+0h䱹�tY���(�Xj�c��ʈ�#���oQY	�������"��}��*����*���Xr@ ��2�3U�B��a�6g3��̟f�
���j�5e�P� h�hb5�.�9-�3E�Ϻͅ*�Z"*ʩ����.$J._yva��;�t�����u�]�Ν��靋��P2o�����3Ao��;;3�j13�`&uc6�	������Ԝ����c��	��9�[P7r�{��/~��
a����,�r�E%�_�Ƞ�J�S�֮�V�B ��n~�5Y�p�`�"���8Qz/�#G�r8zD��Rr���ӗ!
w�ɭ�r8����Je|?���q4�P�n���m�Z�8�/#m[��ɸ�"�^Þ��] ^������:⃃���9hC���8�SHҏ�����FŞ=��� S
�d� ��@�B
_�(���l-{B9�m�۷��`<cˑ�Ju��~R��qMo82Lm�ETm�����    IDAT�� �K%��2 ���I�z >@���R���b�O��"�'�0�ZgQKL(����p�&���:䞩�*j�Y�d�nw�k���r���,��'��2F~8�K3�a����Ŏ�/�,K)��&?���C*NV��|%��Z�m�T��?���A�Ja�(G����r�t�v$���0�-/e6w�=������J����b�ܞ�,���vC��k�x���/����%�kxs���w��x|=�1qe�9�;A�9l��D��$1Y��@0lZ�l�o=�Z���G�:޺l���:��K>Ag�;� �����h�a�ϣe'�F:�Kp%�E<U<��#/����P��m۶��[��ƛd���|�b5>|�\I��d�Uf�Q�"w�O���	jB���A�͐mӖ��N�׸��-86�_w$��%&&���./�/�(��Z�£wa4#�Q� .��g&�0#8�qr�e3�0G0����*u���P%Q�i�;ߑv^�B�f�i�$U��e�.~��fO\֓�W��Rf�j-�r����L&�H����o(�[�K9�@��Z4)�ҡ�s��{�?�Z�n��w'�YWȇ:�O:��6�z��O�A�c`�'Cd��a�WK.���W����hv���Y[p��%7�ou@I�&��f�O��:�G�p��9��0��z� P������a�c�֭ �I{����l��y��$��ʌ�C:��˓�f��<�hfnO��eQ
���!�S�g��J9�d�a�.ʯ)š2�Bah$+8���R��J��rLjD�+�`w/���,�!<�"|��!0�q�jC
4UObd��{|�S�鮖�E�.�{a����z�k�X�b�t�'u������E9*���L-�*S+wz1����w�|o�o�rn2*#C[ȃ|�2Ć�n� ^���>��͋o�<�(x4���rR�Aε�<��Y|�������^t�9�� 6��x�uy3tr^�I�(��@R_|�N5\s���V�i�-y A���5)�� Jnf�6­�(�
2'�&�`F(�
��)����<��W4��~�nobΊE�P�<HGD(��� �� (C��*�jQl���q#��K���t)�z�I�O%�!k>�'��s_�|��\bZ$�#��_�����+�N��ӻ-��������7�D���6����Z6�
\����O���M�DJ3h^�M���iֿDAh��d���$(�x��%q.�JbMj"��#Y*&��L%[D9'��'�q��\��ʥ�'\�s�dGO��b�]��B��0��;_Q��=#r�ȣW�X'<�-���u���x����\-C��X��ռ[����i*4�N��AXԪ&H��}�z��$��<|B� J4�0;������d�́O)MC>�z(̧��[��2"]8
�@ݼ���� H�V��:I+ ��P�\0����+��v��n��hO��2"3E	w�;O]bCP�]�l��DL�T/\s���jey�|.==2��w#�D�u@��?��G��{�� ]���R|��YF�E�m40��t��̺��e_:EM��-��\��Y[}�Rw7|i�y�8y�PJ�mc���W�`.��׊F9�������H��Y��I.��af�s'���=zt���l�������'��B�eՌ�-�cc���N�gg8��rzs�[kL���ͷ�# Z���k���˴Z��=5�D��$NY�|·������1��4����d��&@���l�Q�K��R ��L�ز"�:�dʾ.XH!"�1@��@%�\��f����'s�Z8{����=�
tS���R�#eCus��YI��ܮ:������s��ҙ�������s`ۮzz)U�zФB9�-��g��_���ͧm���^�z�S��}�4Ɨ�_����Uh7]��B.�Ӫ��C�%>����A�%JA
�a�Α(�yk'O{��'����d��<�&GoW(TN�x���}��N;��'0J^d�Ky��<�_�`鏕sY�[�rvu��e~�87?�̏���^������Z+�1]r���q�)Mx���$��Or�B���8_AW�f�OAv&�kƉ$�v�<S�&0u���O�l�mu����h	BK�O؝`�	�漇�|~���{zpq#�F>Qy�է��.U����l�@�"<����R>�u�>��������3ScO/-�z{6c�yy��;����K���O�W�����w��Ŗ����zxX��:Sgw�	3wѓ�eU��<�)V�?fr<����k��M�J�5ԯw���Ї?8u~���G2��}�� �����c'ǣ�̹r8�H+�%B�}<0�xm��᪟:s~hh Db�D"��󹙹���-#�X
���E�j��w楉5V���<����`4���H�!p"�,����S�����m�~�4����ꫯ�1A��6��I�`RJ�X�.�~Z��*��|Eè�l:Bz˾��\y��vU�c��ԝ�+E���(v��w�zy�lػ{���M�(���L���@]�n���B����kZ�,�*V�pc)$���rΎ��B���;���~�}�޺0wx)~���936	���Gb�@�9�}���gñ��_<r�ԑ� V9����\���I=i�Ch�d��ӛ�k5=o����ʓ���-SM� @�T�a��2�V��D�/=RAJ��v!3��f�z��<1HM	�1X)kDԜ֊.j�{jDH 
�J��e =R;3/���T�`�{��dI �89��6$��o�����Ӝ�Fw�h1�j	�6x��G��%�+�P	@��r��uN�U>�%�4��r<�>rO�8á�r���/����+���PS�*.�tHa�?I!���ԇ�N�qA�K53����T7�Q���H]�EO]�EI�X�H�U����_�M�ٱ�ZE��O�L��\� N��f��$2s�M��`p%?5:��:��͖8��pm�P/�_ב���W��\6���>;}�����r�(�@��~�����*�A?73yn��wn۾yt��;�u��O�L
���qG셻qhZw"����Z�D�������?x����̏��e�v��޽�FG�q���Ο<59��y�{>��ϼW��]r����uH��b��q�Ɵ�0��~���24�k�l��K S��~Va�I�|��?q*K)Ԣ����%E��p$Ն&�8�-�r���
��#/j�rr�z,�O�5���>���������[�m&�} R��Uz��"҂$��5�pֹ��c���`���"�y�߃�\ٍ%�<u&����{��E�4���|0�ڱ���ڪ^�If�*�H����}�*
�R$fG˜����,Fn~X��˃ !�m;���})X�:x���|�c�޲v���j�R��5A��o=����s|]����V17cw�9����������׏������w>�(�b~�������ر�|莧�y�?}t)~`�n���z:y߰%r���F^����M��V�A~��y���ԡS�q���0^ �H��&�;�n'M���/D����,3�p����%��� @�\ ��~_�V��/�{��k_���z�F�g��K᜾�#\~C�
Uv=s��R��.��%P/�3�gF�CT�"�g�J��695���/ֲy��l����R�:�L�a"�ݼ�2����%j�9��*W#pp:`&�(5@�@%��b��UU��*U�+�G�U��C�\<�����?}�-�z;��\ӗҋ��yt���Е�hP\�jd1���߿��߻u�??}jz���=`�7�r�0�$"��B[S��^:�J8�U����;q�����\&[��p5�`=u�����û�!�0gV�	�ZT���V�>�l;<u���>Ӈ�f�*�2_�-.)$?�=���E�a	8Y�\�@��흙�~�ɗN���c�#R~W+.�b���)���H�wP�J�c��S.9�t�aM��A�����D#��D<�K.&�˕Ztx;|-%����Х?��%�|�cd�U`�_�`^N�u�d����������I��T����������''���>�Ζ �j6������'���N8�1v�22@) ���j��H��48=-"�^@yt���۶���ϡ���;�ѡ����ƻDP�N�sہ�p�aK�L��_�;��y��-�N�t���C���`I.�<}�<�P�X�\��[0��'`d~�����Q�(@���p�e*�c��.ET�Q��Px�9]B蕪.��b��V�2
"�B���05YA5���J[O�\a{]�-��`e*�M�<h݊�r6N4��c�	��՝�.eZ� �8mH�
��:��q��QC���}eqքu ����an�.�z�(�8O��v��f~s �1d$��聵��a7?�ʼ��$��tq�I���ǧg�9���b�T����{����j%�Ϗ}���~�ã[�B�\�܇0�]W8G��ΣK��	_����6!`��Y���-̽�����n	��:]�5�@�y����Ȟ]�'ξ�8&���tp�7L{��"�,��^h�\,'��.���(!�@��F�E'��#�uD-{&�0��u�A)r��50#Wg���R��&��.s�j ��v�69�a�l���VCA����g���2�k��.�R�h$��гqS[[A�*�=&<*�aJ���_�ڡ]�R`�!pL�b� �=����TZTh�=�N���ҟ�᭍ #i����iF���W8>��M���*�ӧ&���b<����:!�7�E[)�J̖��Ѱ�_���>��n��1�X�	eC W HW��G�U.�d�HT��ʆK	�
d'���`�v�-r���ky\�r�_���S��e8q�q׺
�j*���ò9��b9���ғk;p��I�����p�A<�0Ӛ��E��MY։"/�dA��
���]B�3��/�]��@'�e:ȋMN�4��C��T*��'��V���7�a���߅pi
N�^�(JNZ)�R	7؜UL������Rd�VW�'��ꡈ7��b3�Vsxw{��R��T:�0xӸ݀�v�hQ�#��7�2#V���cF�2_��b���p:?�>z����{��rT�^��!�R6�T��o�e�{�s��~�ˀ.�y�N����"�V��XU���RcŇb�/�PV���[^N!bi�an\�Bt%נ��s��EY��T<���)�Y[��?P*Yg�����&@r{��kZl�+ٻ��t�?�CВ�z��{+OLd�=(E�����K_Q7��U�!4��!J�	Z��
٫$�`/ָ�]R�ɍ$�]��pd�a�#�L��10<D?��l�b2ݨaA���K�Yc�O�@�B�T�*�p��P�k�#�	z��~��d&��)k`��U`�t�F}��Afg�Ca~kF�e���GG��U�*'6����<ʲNO����>�V
B�E��w���?���E�]t
��,�
��o>B�T��(�z�3Rk�8O)�^���([�[9�N���F��ܹ��[ax[�1����Zj���;vm�	f��z�E?j�����s��n�+�G����>�/փ���c�����w{@$v<p�"�w���jݿ���]�s��k3�����E���PM����Uß*��}��#����FO�,��E"���SPj>�yP��}�o��'��2Bެ+�O
ݽ6X����kE! �K�9 �w�/���xc量<s����(24��w�ٛ���	$JQ�p��}Re>my$`�@gbIO�j$Z��Xsc=��E�Ƣ���E|�^��G���)a�0�͠^ճ���V� Ea_ʨ�U�덉�@��Pd̋>�p��d���5��Ӏ�t�ف~ehh7S '.���,�s�zQ�_[��*rG�D�z��A�[fRh��E�@ NF]
�K���ڵe15kI�J�*�e!$��k��*�,g�'�ˉX���Qm};�(���#FZ�6��
� 7���c&Ξ,���+̤�uo�R+�bN�I'���-�����g>����!Bu�d���LZH�_���ˌ���&8^z��8oCUtrr��O������y��玞<�r�����h����l�Sss��z�L�7oe��'�|���  }C=�dr�/~��Q��7�5���N}��	�0
$��,�##.FST��l8r�,���t,�1�O|�w߾54g�h,�=V��&�Kn	�A�n?6,|�������ҳ��,p��77�L��4�02���� �2��Z���[��*���Pa�
��Y����&0C��I��F�W��W�R���Z�`c���H���Z-��r�8~���3����N��4=^��B��?��_����m�nk�����T �M��" ]�����s�?���{�d��?��]�YZJ��gO��kX�a�/�Y�/Mė&G�n�~K(�������S��8�ꁶ��et�fĪ1�H+�^�X�3��}*�:�)�K8r������L�������A�N�E�"�/��X�"ʬT"�m��_C]F{b'� �$#.��n;jm�	�B���f'V�%��f��D��ϋ*U�eU��٩q�[[�U�ڜ��qh '$���W�\�:λd��x�.`)²�k�E��p��ߺ9�Ա�5���"�!�U�:a���믿2��y�����Z��8y�p�x�=_��WC!1��Ú�/��yt�8AX�r�	�ī &�pOmo�g�y��'>�޼y��w�㙧;���Ȩ��V*�}~��={w�3�>6V��o>��+�����aB��P��T׮�;���5f��2=<��bj�-�-��)5�����0�W��NO��*�L=�

DZ��&�JA��U�ㅕr��{��^;77�N� �R¥.dɘ25kQ���	���*�6��m~����,PsB��*؜�5�ܸJe/J \� ���J�^/m`k:W���0}���*�t�I����YT��lʻ�;�3�l}�C\"Ñ�/'�v��G��W�����p���b$���6B��%��~n2�]�GQ?B���`x�Zp9��o��>v�'��^�Ӂ{�,��!$ӻ��3Ο����~z���=T,�b=}����J� ��^*�Ӝp���h����ʤ�ȅ57��[l[yQ9P�B���2.��������)|u��-"�+�%�R�!9�Q$o3�����!4�� �@i�
��0-'�����g�
\����K4�e-כ=����@);�������
�3jb��m����Fϣe��p%��L��L�xz�"#�P�ܯ-�+úgP�fC1_ϥ���������;wt�KEn=<�0����v�*���RV�@U.�-w�e����&E�����O�p���P���{�èxVj	��ds,�m�>�����~��r5��?�%)�!|1v�ME�	�X�z�[��*��|U�i[���~2s��0&%��òF!���C�=��"<˺��'��eU��T���d�W=X��#�y1*��5-Z����3N/#h��K���"B~�l~E��������ZN�]��:�I���6�D;rhti�agU�* �ס:7�&k��:��w�_a;�FY�$��ܗ��y���r��hGp8���a��{���%�[�ٸAl�K�G�'䍬.��	����(KO� V�S��#���_}k�蠽�m�j�M͐��ҹs�WcV��������\W�@��.�"j�.�%�7
�[c)Yڦ��a\��j�A6HU�]e�u���9B��P���9Z6�}(t�ĎF��:�]�F���H����x�W���Hj{N�,��xE� � Q�Yw��Ɩ�[I����[��S��JQȲ�Ɇ$�nj���pm_p����1-�J\�a��xK�R[����+Պ��G���c)���Ȳ�i��t���sTBl�<jr�\����!��iʍ{S���v����������b��W��    IDAT��iT
�.W8�����P:=�ҳǏfЏ�DC�b���D�` ���u�a�f/�lE|��4���l�U����_��L�
�'� ӫi�dhh�r[. !�8nw� O�^�)���в�V}�
�rʰ9���Hԫd�u��ҕ-�o..���ꆑ�=*!'yH4y��^�Ҳ=|�2�*Z���hU>Mn�(i;
D?�U���8�1�X�6����3G���XΞ����L.���l[U��|���Ǖ���S8H�so!�+O���)�L�>3��~9�"��@���Ȏ�/�b%_�`Lb�]���R�Q�`7;�wdQs�$+�^N����d(<`�J����ُCw�P��!|7��N愈�����'�,��c�//D@�5d����Y����W���~J�;�>�a�7�s�	Y���
�T�
�r>ę����aQ'�����dB��c��H���k*C5�Is�f�E��ɷ�U�@ ��'<V��IS�Zt�ER o�j�-�l����g�h��@9�~>$¨'U��ʥ���I٤�'b����y���_��W��B�X\5c>ĵ����0:�4lC�_̂~���Y~�|o��j���߬���;U�U�ʷ�/VD����v_�8�
�P(:8�yvfa||*�F�=�*F#=7;��XŝF��?�b
P-�v����RۏQ=��W��
��c9V��PΡ��=.�s�5�E!$��2�iW',>v}�%��577�����E^X��ݠA##LƱ��lbryn�%�҄03�ht�v0�	a�.�1*ļ�Q���{�&R|4����m�hm97jJ8�P`������Cӣ��'48�
�l.��-��Ç; �v2��,1h��\0h,3QO���4�].`Lvy�01�U�#����t�T���'�֩mMТ\���43��#�G�uQw�H�Ű`�	�j_�� ��ϣ�S�9J�R|�֝���A*(^�G76����|�g�\qTjg�m�2h�ƅQ�,K'�
�겘��NL�S�5]���Ҍ��a�'
_���'}��E��y�!VشE7v���ǟ�������`O��G�-&���[)��r���y`����}��e4$��`���K�պ���*�S�<��L�F`���[��ɤ�K�Y�h	�^�0i�a����u�ёt2�:�.W�m�u��T0�:�͝�S�̐����M�{���W��>�&�C<j(jɎD��&5uw���_6@np��;�!��%��N?�+��q>ԇq8��0�ڹPF�H�xWAHJ�����2�k��������y�_�G�����#��(���i�?����)�������Z�A]Y{l�|_S�̈́�9�C��`L͋S�g<�2S�m��T�'���|��B{ʔ�`m*�U1��8>ZO�ti�����GB��c2���u��v��9�����"z��Q��pBޅ�0k�m���#x��J�;r��F҅�xO�j��%�F����.f�fgM\iF�W"�e��Q_��s��\��������&��G��$r� d3بK1� I�C����� [l��2��/����'#�n���v¥��U9�;e�n[��JD�p�E9��nL�0�F��ďl�Qb�++�
�<X�Ws%4w�B��ՋJi���ˆ�J�x��6)�6ĺ��A���7��Np�S/�<b���Ȏz8���p׃yC��!��uqq#=�Q��d��>7mڴ}$V����ry�{m� M�� $�=��b�Z�:1;3[#�	��%h�m97j���F����B.�0?�W^!�-��>"J�������>U���Wj�7��\��Eh�簉�}	�����s�dBI20IJ^XSbF��Ȏuwr#�%� ڏqx���Z�e�17��[[|�Բ�r6K�]�����E$d妒�T��Kel��?`��~�+���(�R�.Vf���DЧ�A
�K�m۶�}�6Ll��Lğ��᧜[�C<J�����w8Be�ٗ^����.��VJnUҍ��̀-�
u �|!�,��Hi� ��pb͙��ȁ1#���>���ȇX�1���B�]�2�*a2��.��z��j2����s ���2��R��g�,�n!�6]���>�I�!i|L��Xp,���R���6�����}i�֭C������O���ӯ��������H#1��눺��W=mO
�i~C�Ɗ�Kj�F�@5����溦e5�!ǀ����dce�!��U��MI]�p�۲�5���Q�P�\N9��7�!��6�3��<t +����
.�'p%�t)���	�sw9�Q��d�f�X��S�b{#��hQ~t糕T*��_�s�i4׋����Us��n�8�!?�5�`I����3Yu���z궞L6�g��\�ٷ'�Ͼg�Ρm;ި�Ϥӕ�a߻��+���'?}�W��x�d!�q���xi�9}�*v��"$( +�0W"��	�I���C�V��r���IU;Ա�6�u�Er���Z=���l.�r���H!��26�=\�ϵ,�e:^"T:o�&�l4h;�
%O0���Ԋ[��<r���4_O%�sڲ|�qh��
$Z��j^܁L!;�pg���
,Ƨ��ݿ7��ĻL�(/I.��!����9��%ө���0�&ʣ���q��8��)��ѥ�k�N�o��o��S�V����v�[�_dDV�\b��|�7��T�l��uo�-`���W���b.�wsC\��{L��i
H/�0ԣ��R�N%8�	;��W��]�.i�7��A�u\B�pqƃ�-97f�����/~�����?11U(��i�<��޽w|�w���?�����3cF��G��$����(ά���X�Q�:�j\���R�R���p�2pr�r��
��&� ���mY�D�t�`)�|r�+^�dU;p�Q��5?�nj�,���^�$h��zâ[���B��7�8�_�H*�۱s�Ћ
2+��FU6��`	Y >e�;�6��mVpM��5RV9��J��873�H��nX�tIߠ��G(g��O~P�ધ�}����|�g>s�×<}����$�����T.���O��3�{����ѯ��{�ӣ��0l��U�T���݌_-�`�s�:�B�����ĸ�?3�g��?�w�	,��yR���X7��
��� �-����³s��=�J*����8	�-�i�x���9�5�sizbf���㯅�	y~jK_\�j�� /�]��;�7833Cx# J`Fg��^���0X��j��zYQ��5�q��4IV"�^,�2����ɜ^�d�t�u�v]r�#�V�6���j�$��DX�Lm���ʗ�����������c�{���nݳe��׏�b|�I�>�v�}��_~���o�o�}y!	;���fd��=1\�� ��Μ{���*5{4ڇ�7�&���<�p-RnME�ۢ��d���SfR�fxvj8~�q��(N�=.)��� ���6�۱1�ۏ7p��SS��?b��\�E�IDP���g�
�[FF��R�(T?K�	]		c�S6��7KmMi
�r�F$_(q>��6j/�I����S��yt	R�l�C�(^sA�4;m��-���p�q襗'��n�z��{>5<�����K����cϏ���N�~����s�{�Xx�V� ������f�1G�z�/���2�N���5MV#�"_4��^cw�����څ�(�����T!3m�zLΒ�=����2�R�q%�
D���ܐO�ɶ��Y+�gf�\Db��(O��^q�^/�Ю�Tr\;É��bjdd�/�Xk��T��d��G際�5�%�%�j\�8p��Ni�1�⡧F?;ۑΣK4o���Pd�2-^���z��@�{�ܱ٩���=�}�'r@|�8���^��}������������gn.~��y�S�R(�u���.�I�k��A�=FN����Ġz7Z8���%4�r���*_j�#"�Ɓŉw�J�T�^2R�J���L���z���qd
0ٖ�$@��<�:b�man8���z�t�P.��N��w2�\��aU^'��z���, �<�aL�F��X��e��zE0VzH����@��!�����)�K�~���+m�J~���n�c�s��M��{���m9��"T�'�}����Ravf�,7_�z׶�O�?y2�I���`�5����˒h��zә4�n
Rh��W�TqlXB��7�O�p�1v��B�+��-Re�D �Lɺ��nO"<T����qJ�FEL�(�R��a��Ah��+�����#{�>$�P�,��g�+�9"/�tz8��Ė�c-�<G�c74��&���jŀWV-s��L]x�A�G�Z�r�6�:�.M��,Y�I:z<ξ�F$����j~��}���Ʉ�k�t._.���`t��so,�SK���֝��� B�\�w즧5U%-٘�n=y�̢��Q��Js����Ů:75(�����0._h�6W�0v\�A�.p2��Z "�ښ5ڲ�!1����>����/�S_f�L g��	Y8XUG{(��'�?�������v�	�d���@reGݪkz��mi�m��D1,m��^��PD�Yf�u���^?��5,<��z��S�=���
�p��üR,� �^�w�m,���?<$֬��r��6�9�!)��ٳ��_Y�`cg\��<�^9E��ʃ:�4��5�u���U���
;�����5J�^q����g9�S��j����cUa��O��+ԥ!b� 5��=�ؖ�A/�;$O�_*�7ۤR��`V��u[�o���M���GS	4�@%�]��Ź�r!�N`���W���Y@LԊ�JD��1��$�NL���ø��d2�]V#�2�㓦��~�S�g.��fJ���*��)4��r8�^/��No��s:r�U��١�ڪ�:��ѥU��\�c���ԗ{r`��s/'3C�#3���׽���{ �ߋn.E	���ȼ�e_���۶�R��t���P��>�	�慅m���Ǫa�J:2��J��Pac2/:\�y�5k�A�j�84�u/�7�E��+c�%3A���y�w�;�v)잂H�����܂��pm(�������86�E�
���<08��֌��]4�n�7t~F[�]�KF�Q���i�ސ����yt)g�*2�\���d����}�`>�¡�Wr��v:��d^;��ݛ�=�0�g	^ω�^n`0�30\��ffk��Q����4#O��04�dL$��M���Fy�a�6��\d�rǭ��j��t=�P47��7+�~T�S�(5+�}�f��c�T+�KF>WD*�p;�P'�@�S��h��y@f"0,���0��079�h,ɂ\�i��.eIv. �
��JT�e��U.�T1�. Y����2u8zaEu�`;�RdX��p��qL9�S+�⇎����_�9c�쿧\�>������g�#�R/e���jq��g��_}����H��'~}�g����j�P+g�iX�T�D9+��m2\�1V�V�8�Fp����>K���%S���~�"�%cԠ-�Dg��:"�>_0���3�i�Hd*���C�pwww�;����'��v�=�AWB`�"�7y�q^��k�Oo���B������f�4O&��/�m�Xt�����La�X����6#�ƺ�Zw������>s�/؍ڙQ+�-<
O��L6�/.����n��>���?z�7����`8�9Q��pQ�"��]1�:X)�ĕr̈L���N����S�a�S��-��ԅ��*�H�%Hql�`LR�mL��vy&����fWO��H���&�9�G��P��0(f�`��bܾXԂD<������s��>VKҤr����+0,�R>� �i�L�s�l� �i����/3{�ѥp+�nANנ$��b�-t��ķ�����ٵg����e������^�
���b>��?�F��3�艓��������36_�ZI�X�r��f����������n_�l6u1�<����
Ejn� 8~*t(�t��{�Y>_y�h���P�t�Ybo����b�놀�y<>�P`;��*0�E�_[
L0�	J�;q ��:��@�r�|\�`��ҩ�1s!��Q5�p�%��<��<z���j�V¯��1l�|���_|i�������ݣ�Xp4X^^J:���~����n���#�~������ሸ|�����xʴ��"�D� �*����&�[�,��݅�1�j

G�"){hSrs�"]�37����dKa'< 9C �]+���:��G�������d�r�JuS����F�8�sx�O&3�9�;q�e�+A���CԴ;X륪ڭ�Z�/��A�ǋ`]�̓x�!�D�A��u�N�2:�.����B�`p)!޴!a�X����ܾ07����?���>���|�;C8@�9
�>>���}���~��	�Jx��]�'0���.�j^Lv�`�K*�)�e��܀#׷")q�qWȬo�����ZjQ��R)H�J��`*�r��oؤX,	��{������,r��R��<�b�N�%Wb�"��������(�i��\�	Vx��^��D��)�u�]��f!�N�,�JP�|�A�Σ˒P�n,Vʜ^��&��^6\iq�lKD"����y��\/��|�����Q�ݷ4]�:�{��_�*�o2\uO@\n=�tʍ��G��.<��p8],x�á�=�c����O�H�\����S��ds3V�5=�)Rt���2[%��D�4}
@��h�(n����>�ЮE��I��D��q"��`"����V�&K����z{���z�[x�ꦲ��d�y�Q��8=F���[v�9�Ci��`��D�9�y�X��?͸���re"V�Z��u�,��z��U/��f0'���[���D/�T���ea;����G�8��&ytq(� u�HG�J[�C�G�����e.2k�m`OxA.W�f�~Ǉ��]/J(K<�~���H���Je�$�HU�i#�.V�bl���X������ g5�7���#������~����vl��YC���r��G/�m��:�t%�,�9�l7u�o�jwo�<���RW�lY�-/�n	uO9-���.����w��I��'c�\-�^����\t�ñX4�ŻW�a�-�S]斫��wcL�֋v!Ϫ�VT�U�K�77I��i+��`�v��w޹�R� ���Z�]rGK��|�v��_{�5�I��6rB�p�p�z[�jnL�W8q�۳��=\�tu��)���U�G�¦��#t��W��4��y��J{Yix����Ȉǋ���c,�]e|��I�B�� (:��$t��i��`]����
X��_g��j�����,ڣ�Z�0��W���������<J;	D2��\����N`��n'�w"�E���; J��S�]�����S�Y5�f]�*�,p}�����<�D!	��#k)^bT�g3�r%[(a?,�{¡�tV�>:q��t`A+�I�J)���&�r|h:O�#9�,���_ߘ���z�C��J@���]|�:�ۀ/���NWˈ�ATr���R��.3��Ꜿ�����D��z��]�/�.]��*e�:�.��_9��a���5.˘B�%�]nO ���Nɋ1<�s5e�m�9~��6�l��Tˡ�3��Vt�v�|�t��������iF�O���G�X�Ƭ׳m�fR���l^1��2�ڍ�� ����<07��qI�f������v��lt{6���ԪIhw;�.�"rF�'Hleg؁)A�d�^���If�g�܎\<��8xs����6�˹���a��)T�-��j|}u����	+0j7���ϛ�gկ7�n�߯Xvb(E�׈E��x���P0�+��
�R��0UsBl���%.���!-�R㦹���n5>���V�o%�F�g��o��k��6�;����Rɩ��Њ &x�V���-ಣC���\��ˉ��Y��p	��[�PΧ�V��ngo0R�f9���ᒝ+KpﵵE�=g7?�#�Q�~f�q��	�}�۶��#f�k�    IDAT��`��X(�s���E<gI~�Y���(���8�SR�����Y�U�Σ�

�F�a���� >@��R9[�1U�@�fu�]��y��d�*��j����[�J�\=�r�X)��._4>���T�i�B%��rNF ^v-�q��
m͏��F�����u�٢�v�[�Ӣ�K&u��J��U9L�F$����/���uNc�A���*��+�B��{���Z��~d��.�q%Bo01A���@l�]��^b�[槜K|ґ���ת�v�cU�U�U�V�0���e�P�L��[@��8�E�I� �C�4�Ѐ��[D�Նh��"���R-������3�]*�$�+�������s���|4�;pϞ/����^�������g��g^|erv�\��kw���C����{��N��xXt�f��r����0#N_�b؏�8�_���aoec�X��k�b>����` �#,|��7� պ�p'��������+��:{�yti��Z��˪�,ʹƨ"���=�\5�\0jK�G������}}��B�Zź���C�;#}�G9_(%���{��2ʎr���=K+p��]��s��Ϯ��6�#}1��-�3������β�:�/ݗS��<Y3��"�H!�d��6�������������o��cm�q`1&��#���GH3M�3=ӹ_�7���O��7==�D���~3�ﻡnթS�N����n�V�@�^�Q�zCb�!�[Zp�n��鞞����d2.��%�X}y��ق�����Ϲ�@.Q�xt�%(�C2"4�8 a;�#��T�>u�k?��7����#α]�?�/��׿��׿���n��>����NM�g�*���^��*�������ռ�,��y�?�~v�o��t�[��>�絊N!'G|��Soq�A\)����Y���K�߫�o6�8ۊ=�w	�G���:��\�_*����yh��\��T�Cϕ��U=A��D�VDk�'�C�4���^rKV7ͫ.[��Ʒ��F��H8[@Z���k���h޼��n��o����O|}��Q"�{�E��#��s�+�x~B�t�G<C��-v�,��� >l-Ur�n$b���$Őȕ�A=����� ��nu{3�?i��s�J!��1D��^�1��w�,������[��ɉ�w��_{2��KV��u�R�B����}뇱�C�\w�����
S�O���F�0��IN�j��_���Uq��/O+��Z^�uy���Tezܯk7\�����5�6ږD����B��zp���ұmL�R�$>�G�a'�I=PI�0���3�e�jImy����F.��gSG����'�Mq�6��iI��yQ@�$k-3o��ҍ7��"�?�����G�����ݖ��}��P��I���]_ٽ�t2�j���n���O<��a�Kd��i���d�
٥�K���Nť���|��vj�sn{ڭj�x�
���L��m�䒁�S�X�v�������ք��N�H�/
.G�Ü�>��@���K��*��v�罸\��T���=G~>�en�ɥr�ؖXn�0���U���u��xI"�;ڕ����[W�O�Vy5]����u��t���\8�Ɏ��/~񕣣��GN`�ac�4��9��f<w!О��N�-��R������G��]����x1���X8G?Q�t��e�"�uv�X\�s�C.	�v�����hY�I_ϟ\��6&0	$�Д�7��n��hW��.�Ѧ�9�߼rs�֌/^� g�����7��a�DD��	�0��G����e7������T��;߲edd����IV��@_�et� ��d���m;$�q:��}���^���¯N�թ���w��R��TO���/�@*"'l�)�8�:�!S���x�2�&�f�R��+t:�XK_(�u��1��]Z	��Ƽ�w�z��Z�R�����T'�o��M�����Ko �AhK�y�:#jZ�!Ǻ�D�d�-[m<\$G�*�rU)5�*L�c'���]d�J�#�%Zq�-����v��I���䋹Z�0�JD4��X�u�6�P#�f��x"u���'O !����j�i;s&/�E�F�[���E�p�_d�K2��	�Jx��ޣ�
����a�E�E�
q��� �s�4��;��.��=�{���SQ�����s���)�ӛ����|AoP�4_��d:���&G�@ȮT�\�����paR��R�#�?�X2�J�u���=�`e��#ӝ�"��Ȋ?k��I���\_��\xC�UDB}��]=]� �n�>�uC����¬^F�I�C,�#.=��0���f
1]ь��9���s�=�/,?��O�x@����Q��$�ʗK>=L8�r�(�k�p`�pS��>O0��3?z`|�x���P,���u��A�p2���������.�3��<]���[���!�#�"��#]|Io��Ze����')�-!��J�l�0Y?yj�c�$�%sEp�d�?�/(����ٺ��4p��%ČM�����[���4Q�ejO�=�+�C�65�+'O�Y�/Z���1?��Dl��wx�}�
+�w;5���p(�Lw�ٖS╲�g�6LO�`&A��="l��E�lq@�mD���B�z���"���mZ�a&��b��ǟ�(<[��%�x#xȥd�×L��a3}Z,� ���}����}�x��/����w�}x��>��������B��0=<=ur��?0�_~�}�����=��Ï�nX�h,�{Ä�Sn��n
p�۔ ��l���������Ƕ?��w��aN�^'�a��o�cbq	^��$��ް>>44�y�f�+o4؏��]�
��<C��yI��<���O.��F�j�J�/��J�6*M��X�|�����}�;o�zi���#{��ڵ�n�2Mħrc'������ǻ�����~졇�
T�Ռ��w�~T�)Y)��������Js�@8�����Oݥi�ac[��F�]A/��f
�@ 88pC$a?�"X7�o����]@i��.��ୟ��6wy~ߺ �R�\b�&)M0q�^��'&�P�L>���/}��ˮZsɶ��n���k_T�c�Ȏ���e��t��x<���9�o<�ȣGp�d���x%U��5�%B����^�
���52:ܕ��[3��|M�+��9d�csMl`�Ǖh%���}�%��"�E�Z�s�=�lK��s�\vjϒ:v���.�{��m:E>����f�4|�$�D���c����������?�t�[��U�����T(mt�ڤ9���;��|�ɽӭ`�����լ�	{�>�ɥ,��s�Pi��nk��~vW���,;�k�p�TO�z���ɂ�o?���s/�TH�E
'�	�Fnrr��˯��}`ͪd8�TJ�#���q�-@*jS:r�?���w�؁�&�G���\qknZ}M>׾���y�]�o�ɕż�3���v���s��^���N�]����0���t��3�9w�����
n�:}�
��\�w�z����Y՜�lëG�B��G�c"2HE"Mo�Z,~�?9=��7�qõW:�0�� �$�a�s���t���nYNW_�P�>YϞv�zH�����O��X��!@~f?�쇈.�2�N�^/T*V�~]�.�yh�I�����a`E�p�
��`զ�1�
��D�/��m��|B9��K\��*��\z��6�?���G��I��Du��t�5�U��#�݃����=v��"o��u���|�l<��?��R�����S�\������Z��Zn}+�*����}��p<F�Z)�!+��0���eA!�.gȥ.ir��!>��G쇸�����N�����r@���B(�3���n� �b3J$�˙% �R��؜��dz�������Z�ۅ�'�����.VJ�C�&*�X����Lg����c����ݵ�����mV��ʯ��lÆI�Q��Å��[��i*_������[��S�!]&Tn��g����Z.�b*��������O.�-e��W����O\$��u?g����z z`����{5��i��v��`(��v��1�ehk:9x5KB���?�����\�Z&�L�ݬ���QaYD����%ޑ1��r239�Z2/a-;���o�ʛK� �A�3�Rt��LǺ�䒷\j��хn,?�ʨ��E�Cg�V�h���W#�@��}�Q-���d ��EO(
���|jfK�t:D�H��a��Zs�p,�Ǖk�'�/�{���Zhl����D�	��r����93�zI�Q����O����"L8Mv��(r��%}z��e� #�F�b�{���8��r��ю7.�$�	�D3tZ	�y��WOZpjl'�P�It���e��������N�91�7�&|���L�L�)I�a��J��L�F"���B�@{��$�=�����&"�r=��&q�옣'�I��OW�%�\�rIa��I#WXI �W�<��e|��'e�5/����[~r�v��y@R7e�P8���g�T.�`4��y�eu��D��x*n��iJ�_/�����M����'g�2�Z0+W_����4��##�s9۱�Uß�n� �w���%I:�o2Q�+G�D��ǹ����[J�������sO�>|��E^9r鮷��]r]oz@2����n��u�����īn�L_��
y�����U=4�����Xlh��{Nwe���n�鵚!_,Xk�ysң׉�D��d�3)�|��P�	{'WNz�Ӭ6�\��w�]yμ�g�����N��t}9�(u0|V�I����wz�܏^螺_�c]�xש\�����d,I8�S�F0�h�sD��8�Ғ�4�7m8L�\�L[Kė$�����������<�Ю��n�ʹ :�+n���l˭p�����3��Y��gx�1�lT�cZA�9�Ǥ���R�]���IHTr	y)�8�UPlj`�dO`ۦ_V@���I�E��9w1�<rٹvYJ�br��؞�N�"bx��Qm�}r�fej�i-
��t�Gī�Z�Tӣ�t��e($�u8L�:BQ��_���<������}��C>9>~��A<(���Hyj��"���Y�X�+����)'H��������y��Ձ�'����Ԗܯ(�:@ݍj$�MZ��/����T)W�fXk���]M���F���H*�aS�CѠ�a��4�*�$�D |��N�r��r��S{:տ��;��l]oY>0@��f�$j�c����kբ���/��>����k02��>��\�A�r�%z�����g�O.E.A��t6�*�eL�ȏ��NhZe�7��J\�����N�Ip�S���9595��kɮt�k 7Z.�D�	��>[[����J�ez׮�|ѵ�^�V�����Z��:������@1%��]�X�9�$�x~�f��?�\��L�����H�OO8l���@�D��|۪��{w����������N5�ǫ���ß��W���R�j�Xҵ`���@�?�G+�W �t0��fź�u7��߳vm� 0�0�1-W�����!Gs��}h�-�ͯ}��Dv�z*�3P�e��tm]����� ����t�E��(�EC�	o�Z�6Mc�E�_׫�x�V�oD�N>|�a�x2�w�57�]�����'?���S$�>U��$y=�a"�_!�ˌAK�\wz��&,��jO��Lb|I���az+E��>]Az�6⥓��U����M"�e<N����r�`a<���RBk�V�Ɗ��)�c ��z�q�5�?��o���7j���{��7�>=r
YȻz��WW*W]w�{��&�Y_�����"A	I�hy}f��|���<��ܱ�6�=�->p�i�-���+�z��T��<���k�ך̦5�:��gGd�d���J�Ń����W�1��0-8����z�q�m������z�_z�b��r�D[�Uũ��Ç����6o��w������GF*塹~,4	G�+�緥z'rىk�����c�GG�̺y���Hh��cT�E1��&8��y͆�4��p�H�s����]�+�%�(��]�����'���ޕ@\B�F��;F�}s�n�'�E�T�6U���ʯ����V*G��'�ڹ�ʫ.���|$��h!۩L7����K_��[���������'�:tj�D8�751	�jԭ����q�qR9!��
Sa>�9�g..������ډ,�!9�*w�λ��?;���'���N�\�렄R ��
�X��:�ȋ7nZ=�i4r���\�I�����C��ވD�����㤠��٠���n����r�m���.��
w���#��3o��x�rjs�G��%�l��%�����'��:���K��:TC9�a��F�eU�\���6�]n�إ7/�vˍ���d���zoHcp����ի%˜�����/���>u�X0z ��o�|�}ҩ1+�a!�Γ��o�Y�n],���E���E�e�G�#���&����Ĺ�p�$�@7�����ݘ/T���xq�/Ыϵ��ƑAh��yP��'�XG"�Į��E�ĺ�%�Z��eە�ֆ[���DCk�/���t�����HK|��i�І�W�<uǙ>������Z}�e���;�0�Z�P�]��Y��"�sml�c
�����W~�^i#F���d�J#�әN��TF�Ѵ������ �(I�Z�1!b�nPL*Q
c5�`/���{�<��W�s�g��>k��XJ9C.ϣ%�\�+Go�]aBD��p�61����.<��N��ǹ˷��53�E*zT7�v�J8�'7]|����ٿ3_����%�@���FY���*$se�ss��ʅ���!���������ݛ	�(���K��b�L�)v�nH`��>o�s׮]0��T
�X�	^=P��䕺�m�R�Щ�M@���'�͙\zX����p�4�e������ݟ�4�Mͮ'� ��Ih��F���aMKy�ˀ�j�X*�#�H�Z�h����"w��1[yr1pi����'��|����=�_4�j�epϰz0^�Vjf �����x��nڴ	��fنß`t��s��e�a����󀀐��K�B�d�-?���mʖH<�5�|'8.B8��,���X��9r��Tn�	���خ[= kI/BhnZ��cF��F���t�'J`���8�,]v{�����>ǟ�N����\b�9%g����x�4	y�z����LCH%"u�����{uI)�����s�\.Z���]��#�H���̳�'���)�����$� ����S'n�拆��Z�<���\q��[��J���Lj��{�~��.�ҳz���|G�:rh����ɮ��4O)j9CYVHLG�X�1.�s/L��m���_v�K��-�$e�v�����B}-r�1\_��t	%t�LtA�"r��s��O;��ܶ��Z�?O<�����ҧB��mc�C`�$���}�SW%�u�>	��ğx��]O���[׬^W>�{�큤��K̃�u�2�b�G^rï^t��}{N?�����D���(�5���0�g�� ��?����y�A��f�v�՗�ƻ~uӦեB>���S�Ѝ�-S��C���}������!h(S�L|{Еc�93���6��{c^���}��|����gHlYg�Ȣ ���2nd����-���ŚA\�H�� 迓����vox���v�U�n�S����?�Iױ�P��Ԓ��~����4'����>6��ٰ�"��f5p�vã�:`kvM��tO�N�u|4$a��ob|*OG�1�̞�r𻎰*�a?T�WAV��>O+��*�E�;$�K�I�K�!vl�#�Gʕ��H�P/3u���G�@��T��Ȯ��4[�F��)�E�ڲE@�@W,��&G��IR���&�lym�Գ�BR$��S�ZIU���XN�����|��UΕ͌BbJ!m��>����6�������ʀLc����&�1��g��3����2�g��/�hUg~%ڙ$��\    IDAT�D���f����!=}�w�fNB����i��Z��K�]]��(c��ѺD�|Q���&�#�/0=ݳ{�n�.���W���V��S��sO�K)���t��w��͟ǳ����6�XlGf�� Uw�AN8�i 	H.Ȧ���?s�p�ȟ����׏����VS�1���ɇw!G���UN��f�m�INژz��n<�cS&�4��� ��ZXk����_���U��7�۲�ʧ�|4����>�_3�~�\�~h�ڍ��#��?|�ѝ�7D6�#ÇJu-��5p�>qш���x�
31��h76�^���`1�	6�S��q6R&���R)��Et�1�w8qi%�B�d�T
�6��!�7,O~z<F!�	)�H����ԍ�x.<���XnB�n���0�L��a�#�1�����	WrnU_ψ�GQ'��e��*E����4���C��d�R��a�sP���@;���$C��]�$l�O�F�\�s�)���A5�K� ���ru�E�Fs��ó5.�/�c8K�$���z1 5��B8�*�
.!l�C+�dQ�A1�PL��h{:��TH���<�S�U��~�xSp�w��1�0i�}�U�O��y\����S��q̦�	F������2su���]~r�Ry�!a*$T�b{�I͉����}�;���ӿ���t�����U��1����T�nٙ�՚�G?�����Ï��ĚH4j#���?C3�VC�&����� 9�cّP���¡@K뺿�j���	J�	��4
 �8qS3Q�S��LL����k)�iY5Ǩ��~�W�����Y!O��5Um�vr��K�5�Bs6�~���`d�d������,q͖Df܄"xL�P�0���R�Kǰ��B)Q7tL�D���z��S\&8L�)��}pN������\Rϋ����J*.@�&M��(��g_?���3�g���g*����=��EQ̹��������i��[�W}�F3$���xN�TQ�^���^�����/9<]�+��z>+.�&;7	�'�_�f����~p�}oz�ׁ�M��D%W(���Lq��"�-ԑÅ �2�1�TsPx�K/�G��hOW~�y�j�������F��s6� ���l��ݻ�S������]�_,������I&�-N4�!̊4�l`�h2��MO�RC�N������$��%��+�e��6���gpP6	r)VnK^il��!�^y��/������f�Vbo��B�>��"	�F�����W�4n~^�*$^�n�8$�ac�����Z�H� ���EFø�ȣ�,:��r<3����Z�B@>(,� �	gp��;�=B�f��m�g�_�{�����Y�O����I�y��?�
MN_G�l�������K��3��`��:�	�0�vK���`�ĥXA2�d-��VD�/a3�`���g�-}a>>g��A&�Y�������sa�ȥ�K��V<�*O�s����u�6�2ЖY'����q�1�^!�����'��FG�=�e75��Bj�i�j���5�n��b��ǳF�G�:�i�gئ]'�O'��;O��q,�(K�"V���r�e��}{�Ӱp.L$�Y�m�cj�p�;?q|_yz�H���!8�y�(dU�Pq��R�)�2�h�l����*sAB'>�R�Oӕ)�g����2��D��;���o�<`�:Y6�p���X~�:�Nh�l�\!GV7�F��,�#��#�Jb�f��E��V��N�(�"l�ee� ��_�!������\�ǹ���Lu�t�>��nsF��>������38k���L����L7fReyS4�}u1'�5%��.��3]H�<Ӿ�m#� wɱ�H�ۄx���d�v�.�z�t"�.����p\]�tz~�G!/�XAׅ��h,{0��c{R�����������/�$�O��^5t�\���ҽ�N��g�@.!a`3<��!*5��`a]��`WD��x �)d͇{������Nwf�Q�xٛ����z��Ѭ�Qo� ��������zi�����vgc%�u:�n9��`I	�y%T�M��xè�xV��\�נ�5��P������z��l}H�f�UM~/B�T4Y.(�V�T����O���U*n�b�D�4%9������<�a$m˄\Yf�)����i�>�y:o�W���#&�B���p�9԰Ħva֐.���_m�-�g�ia�h���k�HKڅ�R� �k�_ܱ�"ӛU]�Up�|Q�v�Q�����W��}�:S��T=SXK�@i������h����ݙ�^=�n�MVa�U-M��E���w��FX�c0���˕pD���O-u9Y�������<���M87ٲ��x=��c{���A�я��U��qgfZ>m��(+j��%{Ŵ*4�����64_�Lyu�a5jF˫��ޠmXZpM��	�<���h|^'���p�ܰ[�(<�d��0�.�?��;��b�N�g�K˶���-���5���>4��gh��~�F��� 5�$,��5Tu5�\B6��®X�0��r$'��ꮖ����Uñ\��>92��o|k���ɛQ��kB~����x���0��U���4e?�:��@��i����Ɋ۶���J!�sȥ�ԑ�Ș;�V �5���, �22�2'm����n�4^V6���Kq����B�f�n)rJ�B`�0Y�%��9�(���"@�����ԋ�%��!p�勏M�k&@�*k�Wg%a��fz0\�����8�Pb�8�ܓ%}w�a�Z���("���E+�{�K���0��f����L��C~_:��[�'�6p���K�i>��|�ӄ��mիf��L���)�I�1j'�=9:��^��R$"�E&&&׬_u���J-Ȧ�:�< 	'�$�
*����ȟ�c9���5j��}���V��h��9GT�_���ݝ�?�ѝ�j�J��s�e{;ͼT�G���dx��ã�]?�n��ձ_�%�:�d����:� ��l�i6l��h�[VQk�%"����U�K�O���y����ń�pn|�-4�e]�����߯��p"�PA�qV�G�wnE�h���%!ͼ'�J�΋<F^뜅�L���G%�*!�nj<[��~ȸ�V��X�_�'n��G'��G�N��켳�֍�POP�I����)t�Z�-��L�SgZ����<�s�@�Ŏ�e�y]�e|2��1֩�Љ��~���rٿ�������FP��ƫ�Q���M�*�����BG�fH��dO�E��r��G7�����t͙X�6��2�X2���-��5�Z<'�u���c3�'RCXEx�J쉐�'S��8��B���_��44b]W+ڣ��:q��7�G��P0f��c6��Hȴ�H$
��h��0j�O�鳻�ؘ��*W��)�n5C�HK�X�#y �/�����ҡ�/�5� S�Ee�f2�,�I5[\ٳ��U�b8��H�I�&2 K�fJ�D����e�u�Wa�\��Mض`�D9���>��R'H�7o5�;���:,�4^r�aw�%�t�cц����@&��ܱ<�-%����,L�0�}A�Rn��0�ش��d>.���۸-Vke��KQ�s9MNy�� �[�9%��J�h}��X�gE�V+F$��٦�����0á`"�������6���{zz�1!�Uc8 ��.��rճ�//��r���X�K��\�k����Qd��~Id�`D�X�G�ݡp`pp��O~�{��A�/��G�3�.F~�g�'��9s�|���[��q����):�I,�� A��݈�G��@+�!-���P��4*�aփA,K%��S�z�{�'�L��)��iCJ^�Uģ"��L�}F ��#����ͯ~�S���c�N�6�AY/�q&��k�F]�XĒ]$��l'��:��U�M0���()|�r���HB?��J9��L:������?F��T&9�����j�h�9P����%�7����Ǜ�&�ih��:����|��E��[BmU�bMW�?�O�fW2�u�6;<�he2"�Xؒ���i�lh� ��Ӵ�(JɮX8T��/�1����*b�͌����X?x)��峎3}\D�s��J�a�QE^�zh�Z��)��yYi�{�5�Ӷo�<1������3�󣉳�Z�4iW'�!#�h�xD���5��Py�A�ߌ��R	��zX����y��d�'_����������n��rl-+`���X8�?1Q��w�Fjz����e��I�q�H1�b��y�Kق�?QɈ/��p�+���X$ĳ�r@|#�FFp�)�D��%�5�^�d�kdT	��<�`�HeA�dNia�O#ȥx_0YdZ���f��
��9�i�Njd|��c0S�촰�ԦG�m��fA.vÈ���(��N>�hZ�iԽ]�h�ר�U��Qo(���0<��rR�9���	�Y�{�	dE&�P=w��d�H(5�MK�%7�z����֭�?��g?���;�@Foe�#��@ ��X�d����ғ3o�I
L�:u���[_}������K?����u�c�w���P�F��ض�:���$1B4���Jj9$
����e6y֨�3]i �T�����o�uC�l�E�3mq����K�����Q����~�TB�]M�����B����ƕ�5f�A��{�1;u<�^}���}m&�E�Q�x�x@�|
����j�������i�+�d@y^��u��,se	�-�Qef�E"FQ|f;�y4���aX����]w���cG>���#��o��o�*ޫ	G "�}f��[�h�/@v����S�	?ah�T�J����I`ò� N�d�
��d�0%e��}a�m4�)�ݴf4!�07��	��C��0.��5m �YF�c�d�f�"Bu��.T�Z��yQ#ȯ�F�\��Q�i5��6�@Y\ܼ-�,��T�@V�1⽳�4ؼWD� �X���C�RE���J�,�i3�E��G��kW�N�+[�2i���PܖK��Qb�~�/t�8o�]����m��~?{̭[�"^��^�N2Q �_C�\y�ຠ������z4��Za|Z�6�-0 ��<��A��H��S���ډ�X&L}i4�U�Rް�:k���9+_JB1�̍���~����Z�[��%�{��`�K��Dp!F�@�n����_��WO�8����u9�m�
ǹծ�/�ȥ;X���isg�����/�+J!{0I�Ǵ��PO�j��&����?O�G�a�"
0��G1��\�f�<v�]�8�	]N4;ұQ!�Z�|v�V��N�L&b�|������ޝY�j5�d8�=u&:��+>H��C�q@i,DS�ݘ)���4��}�2�>�#>?9�1���˿|ۦMCG���׾9=u�TW-ô���8��Y�H"����q��7�E��u���A�jE{{��izR�.�sq����Rf/�S$]N0*��
����AN�zr������^8�k��@/�FA�)�N�R��a>��"���"��X��=�5��߽�{��޴��P�;z��0�E�:A�b�,��5IWi:�C+g2��Ng'�����'�}�����%!i�"�޾rv�-;����#��4Bdނ���T_�j�D���W �.�Ӡ�
�y�D�c��a6/�\qzr*�?�Gq �D��U:�.O��bB�t��"�K�#2�Q��Уy�~a�\*9P�
 ܱ�A\�j�'�SL�I��*.��N�}�-�J��~��@����w�1���gZϙ��T���=�B��#����c�`@/�r�Ұ����(m7ݲq�@Z�d>�;|8}����G&��G-z}kz�Q���f�Qf�#c��~[U��,�j����V��aֈ���7����y�р�;et���|��n{��W�ڹ�~06zȴ ��6�24Sk�th��~�u/��_yW�d������&��0Z�J�1kߐ��Z��W5��'�K�ܫ�z�9��A��>�waNi��%�;&s�F]���25 �EE�P���ݪ0^4L��Ⴧ��$$�xQ���R��z3�>�Ah$_�^!��c�N�j�baz��/�N]o������@+&����Y3����$���Y���7��7<��Q/�{��eONg�KW�)p?[�*r[p��"����?j��~��h��f٥����m�m������*8M�O�m��!��{�,K%�K�H�h� G���dQ�z�P��F���׳! �͡���!���ȇ��(��P �<���\���6ۼZQ���Q���e+�k4j�@�%�����eh���K+A?�e\-2z`}.���O�஧�~�R��KYȜr�?d±�d�'��+��2%a	����37=0j�Rv@f�@,� 3G��N��9/�Z!���P/1�=&��|�vIN��;y��S;w��F$�$DH�P��?���f2={8]�W�lOWN�3����Ž�p��,��.ڬ`[��=����z���3�ϝ��8v��C\V������h$R�	���@V,��-[������ �s;�jI�M����׽��W^%�ѭsY]�r�
N-]�	�⿿0���>t3�|T�.&������G���Oe�2H�(w(������Ӿ8���Ŵ�7�Qſx�@X�|1KĽ��jy�;�0��S��`r���zs��R� p�W�ӂϜ�E�FO@�w`L�@lj�n.W+�H�)�J�*�N}��E���OX�Y�;�u'0__�ϷY�{���ǡ.��hw�갯q�F�/��;o�{~���ĩ�"2��&�<���.�r��W_3����H�\�kXY�M�ĊX�$J�V�]���P:4,�����E�YȖ���`8�m��V���b6;��>"TR�lT�".0�������CZJ�醊e�ؖ�@��a����t�|�q�{R�V("��R���+	��ӕr�n6�WB�b)����!.�T[	U�"h%��c낽=μ/��!J	��1���Z٣B߱��SH�mQL��G�"�r̗�T�����?�V��i�Ѩ�iY����wUsgZ�,X:p���ۇ��Gnx�U������?�����7R�M@1�+?��;�#��5�d*�~4��Ll50��݆D����@�Ny)� ����_Izq.��������ʯ�����iF�
��G�L,Ax,+e#��h�H406q�c�+ì��?�y�E2�b�. �����ډ�v h�t��ۗmؓZ(��7oN�}/��w]jd�rx����Uo+Ҳ��}O~�꫟غm��n���?|�����>6��g�ʕ\�q�f�b��8��@oP�i6�1=j���f�A��`׬�-��"�F=���i����sYC��1L+�>��h{��k3�� F���s�֭"L֬� O$�OOjv=�N��j�K����14$���,�~B1�W�ad�$�Z6U�,V�Wl}����Q�Y+�{�1]�t�A�NE��>Z��\�##��"Ԗ���F�V0	�6��������w��}�O�~rס���F�G�a(� �(�D�}�F�l�\��5^OupU�m�I��6�ߖ�/kj�	� ���F�8
��X�q��%�s�Ԩ���b��d��=22Ft�d<����`]mv��u�%��K_|����N�)L�B�x8`}l5ekp�b����+TD�{����8$��믻4�d*o���ދ&��`��6C�
�%�7z�X
)��(���"�B�ث���%���Ɲ�󚱼?I�� ���W:}E�,�t��A�s����k�B����CȮ��DUz�Sj��[A�?�����a�]��/��@��3����j#Na�Q��"�6��ц��J��aL�#��j�Z�ɏ������E�N2��t|�Y~�R,{�)"e/��0��Y�X�Q����W��57b���#����ɉ��/[�j�Ԏ��=26>��^v�moy�ٲ����)�2��a�D��-�(���h�JɎ�@e�$���    IDAT���R(�	�b0J�`�;�bH�2�~T0�*��5F
oJL}�!�`�LD����I�	۪�����
&�Z�D���R�^��}i͓�q�2�@� 2@Ϳ�ܶ���}qOF;}r�;��棞G�+�>�<�T�WS��0#e�����M7��;��"�>�����Ŗs��ɮ�قO��B������^"�uwezz��a�Ph�ͧ>���~Of^q��S�cGG>�+� �[�v���6o�R-���݋Ƌ�6��<��{����v��k�nݺ5ED�B�Z�"���C�yϯ]y�EA�+m���N&�%��Ii�:&���T0��E��C��bf��!:��!�NN���-!;9�6�
:@\"��E
J���j.-�?W.��md�)1+s)\?�z>��m�'ؑ,�(���"���%�r饴M�4�� d�9c �z���011�f��&��2q!���x�<Y�U���4��^�v]��D�ǶF�Y3�=��CO�ꎫ��� �J���O��"�n�	����[���M��v����=�ǧ�[.��տ������HR�������(��x�p�e���#?|
�A�Z3i��
-f��b+�D�P�T"�J]FwwW�@W�X��p���+�oW�M��U�&d6�H�z4��Їm�9���+JJs�Y��!�L�Y��z}:!1X"al�q�a�1�Y�0!�j:)������Fwwxj�8�8"��ނ��S��{�n�>/Wa����q�#G������v���ӓ5�
�����/U��)]��8�%�A4м�X"���S��wϞ}{c��σkN\b��.����O���	H0d�]�]V��L��-�0j�(G�J$�r��t��cG�_��[_t�E��l��b9<[4
J���k���Hd�ݳ�ȟ��_��&�A|�0#�3��>D-���_���Q���aY�Z�7���;�J^�q��ڂ.�5K����\��� ���
��D��YG%��3Bu$ȡ"��<1u�X�2/��>��N�Y%�QW8Q�#���&O�4f�<���!�t'	����x��X,V�9�jcllƚ^bs������"�H�+$Y�we~Zt.�yi����3���X�[׭���]����c�=}�n}��Z�m�Y��**�������=�=�ӧ��p"���UG�f�>~�zо���H9BGܣpV�h6cAb�[Z�Z���`�Z���j�V9�bq}� �=$���{���A/��	��b��r�X5�(��x��l�+Ӿ���3~٣5���gS9+�] l�i&�]���]��#����u�E�6]���c2J*u�z �r!pi���X4Ƅ�>�f�V�����0M�͞X<MĦ�vKpU�_�+�u�d9�&1��	X��ʁ�G	�D����Ox<���$�5b�������_��!��ɮ�6[v����,6
��E�鑑S#�:VO��3#�)�UfT}g][�o*�59y�K_��c��)�O�|s]f-S�SCo�W�X�n޺D\����/R�Z�=@�O$�b�,*"��\�#�gh!3:|��4 RWsY�HQ�٣��,�(��]�Q�����f��&��c&H)���k�?�D�Ha�!?���+����U!5�Ù������(�%�c�~�jժ��~�T�j���rȥ�}�1v��Ź�;C�K/�0�O��GJ���ZkS���G��2�v0F���o��F�G��t���p�֓ǳ��NL��H�^�I�R�٣�)�;-ķ���ܹ�������{�P��>u�@���4��o~�F��b����ۇ�h��qB�Oe�z����?����|T4i�d�|�1�@�w_/M������M�s&R��,`e}c�	s���|��]+����5=�f�qQ&���:SA�lYN،�3�lA$�G���( �*�h,O��E�Q�\NJ����5�e9���M� ���#��C܉)�Y�{#�f�gr�%W^z�@�<��496�y\�u��`��z8�җl��%/é��wl������ @��!1v�h�<�)��h8b"�9�ۏ-|"a�P4�ۻ���{3Z��</<��u�K����>$����%B�z��E�#|�j��s6]e�^X���UV<�>�xő��X��\��;�y֍9p>�z�˳�w��x���Ay��D�}����,�I��8����@��	M�Q��o��>6|��Cf3��?��K�>�=��a��d�H����F} �tl|��gw�B�]�"<3:5w��=��&Ih�=FI�+F��47�\���T=Ѵ�[�n�.�x��!��@��z�?M�m
G���,��]=@\O��%�93{�B2��L��m7�@��s�r����V@J2�jF��Z���:����X�]�~l�L1{�h9/!�Y�FǊNs����4I�c���uG�P%��R���|w)�;�x�p$�\0�5�-�a���8�̲��>��ˌ�� ��F!W���ǲՏ��H�@1B�tTDqI�\5}�u�u��N�2=���ِ��+�����w�s���r�_����4[�*�c��چ@�#�k�����}
�/~yM._{����i�t"�WW��;0�{���Cв%�:�h*VPp	ì�OLm۶���� d,(�K�H<_ �7�7rn\0�2E[{��)���$I����=8$�d@"	Û,"�b��O�psq�Bݝ���_�T=m��s`Ac�R��Ž%��_Q~���"���PK�(K]���?�֧aa؀�Y}�Z1��ky�L>of������S�L�x2� �MT 6���طP��Ꮠ���C�x�e��Dxp�&�)��~�i��r65cl�8U-��D�%��V�����-�|Q-��	Pa�`�^a�A��0�≨bĨ{���*�.:N�N�_��n�nt�7�V�:~rdm��LW
�x,42|
� �-B]��8m`6�2�DP����{�V/gs���;S���f�8	o����֟�gǖ���ΚmN���&U�E�:Ar-N.�t����q�����Ya�E&�I��}Iͷ�_��7�D&#���a�믻���"�ǋS�B!k�ƄM,���H*��'��l�u�Ҫ�o��J�Ox��A�����R6�/J���F�(�xg	����r��i�zDXI��&٩�c��ކ���^��h�=H3E}z
3�p!���R�m֌r>۲m�Ƶ�z��"j,���
-��	w�U3v"-g���݋�8/�3h��(�}�߄\r;����jV�<0����-�KA0��*�p�522�0:i�~�M:ݞCguI��,�.�9��BC�!�|E,c���Ik�)���
���hBi�K���,�N�pp��7���#��o��o`���I|0�����l�RG<,��|�⢽���bً*�ٵ��a19#ͭ(ʽ9\�+�q!@�|>�=�?t�'��a+�ޛ޷�\+OL���}R�>�3���b�����6%��^4�'O���ޖ�����׿��
�*6e*�NJ��! �M �����}0����+_��`�y���Hֱ)�Ɉ�P�8��ܪ���e��5$��O���߱zuω#��N���c4>�Dg��A�-`ǜ_�W��/
4y��	�No�������&�ڽ���������W���Bxmȷ;�]:.|+[�f*��D�L&EY��I��r�Q+�}cc�w=�o��c���+b���T��Ԗ�K8�NOO�������
<emO�P�%D�kE�{jf�׌%���C���`,f�>�555������Ɩ�dEu��cP�8�Q�Y�>*�q_�,�-�Ǆ�80�ت��J���s`�-.�<{.�@r!� 7���:]����"Dv[v���K�
����lde�ㄍlUlW���LM�d��|��~���۞�y�/?��/}�;djX�f3��1waN��T^>�h����ƂPZ~r��B	�ǆ�^��d&�h�G�?�淾e��˵	�Z-=��+�]3��W"xe�J0�ٷ����^|��Ȍ�nY�c����@��ff�Ee���C�XZ�C"����e�����`��CaƤǀk�=��Go�h���"1�L4j��\����!#����CA�	�I6�d��V�i�v�䓀|�A�(��?'��Z ���Sh*FQ�W������ņ��&����G�DR;�R1��c����C{SD#1�Y�� ��A����b�F�	S
V����7�
�l�R,��)� ����oT(f�,@Lz�6���c`h��ќ�{$N��eW{z��Z�#C�5	�1�*�� &����X�x��
'P�x�R]_vz�7��Q���"H�*�Q�>ڽ����
���W2!���a��G�H�Z<��'O�<B��\����#�vޕs��{E�zv�]1�P�)���DK	�{�΂��-��Bh,t��K����]�^�f˅,���׆I�X$�<���#p o��$2�Dy�:�m�����*y7>��o|ë���֮z��-[/��1w.��b��>|̯��Q��NWw�^�v�V�3���;��"(���.�U�D'����/�W����ʞ���]q�k��l߳����G7]u�t�t��;cçw#-���^6~�t�������0՝��J£2rh���ꆻ�j-K\�0z�$���o��m_5�Z�v-kC�`<��V�J[wL/{����l���R��Ӛ���Ţ��z�DN��H'�xdx�X�8uц�Wl����Pg�P�S�̣ pZ~���_���Px�8���+�/�]���YEf���<�DčS�����u�]'O�"]�$rd��q	a�ĩ6M�1-�i��HQGw��-����*q���;�;�Xd�V��R{�<�O�lUz;� �m��f�2}��7�gU	��Qj�!��g�V���� �%!�0Ք��ݎ�&��\0���fC�@	�:-�rӠ��q��	���zM"�ƀl�Bcܟ�c���:���$�w�M��m�ʗRܥt�7�rA¸E�\[���ޛo�� U�Q٩��S.�U2w�v�}!�̽ڦ�s/Μ��`�'�Fd��sh�0�t��1�� # ��c8`k�s�Poϱ�H�5}��7���?��+��\(���f�N����$�Eg�������M�^+���>ł,��E�,�Ǐ���:璭laQ��$dw�� R��c���_�ˬ��W��_ݿ�������O��}\w�@ �jX�`���\~勴V��;�?��#����1b7FS-{�'R`(cO��Dԗ�db1���ݻ�_��O7ӵa�L�V���+���O9||݆ͫW���F�jͬ��D
�*��f}|���&�GB���u3}��pp��'��n��zׯ�����l�;EY����rM�7#}�d����J������h�ڣ��J\��P��\�VB1��)�{<h0�O�iMĎ=�0��h"r��Wſ�g��	eFK����5=OEM	</!뫄��iN�C������[�nM�R�g{�r�b!s�q7'Υ�}Y�#'��by�iT���j�J~���)�	�|Z�D�5[�)�qk	��g�E��h��;��S�GV�a���|H���5�bd�>5��]�ʳ^H's�\2zz�j��S�\�%񌡉"Ǹ���nU@;9/&�]�nF�[BL	���r
�PQ����*��1�IDxZ����\�#��D�E{̷�F�w�cD�F���4�pc8���X�8]/�e|[����_����kI,�!�����~�����&�z��S'��s��@3�B�H�
�H����̰��h1�������Հ������${.aU|�=��}�{����m�p�U��cwﻛ���$T����/��'��Ԓ��`�?}��>�x�l�kI��C_�읙?j8��'&��`
�92��/|��_�:���t��'���A�����_e���x|{8��$
Ŋl��\kA&ȯ��af�U���w����Q����c�X׭�܀!�H.�7��B,�b*�#�	�uLX�-�b`�]�vj~�5M�����q2f�3U1��X�5�����_LV�j���6	��%���kOtI榖�N�|x������j�����,�x��1�ҳ1��$۲h@*�s����;j��`gy�z�~[V���F����%����#�@��#��)ʉ�p	E��f,��'���@�t�aC��f�E��D�Gf�q��h�	��%��X�QN����?q�2��.�m���{���j�[d@qU�ɀ�-�D`ѳdq�s�J\�U-LD�L'� ���C�<N:qV�t�!pb�����i�
�a�t�X����a���0M���<A2D�oz���/ }G����}�ӟ��SO�fFc�z���C�lif�n
f��Q]a���P�����s��H�ǌ%�$긬�MO�g�4Vٽ��w����zѶ�[�����!��^o��]��k��J}�OG����{��x4\������<;3u��3��4�E+Uю50Ud��g�����tuخZ�ư�h�ر�^��W��8�J�S�v�������#�Ø5}D�I�
������g)* ����_��0!�`�X"�A6փ[��c�5��� (���(m$WȒHZ��˨�9�ۈ	�S����+!2Ws����:��[��!�@E��ʎ�%)&��H]��5�{��+�Y��"��9�삲�il��{����=v���ٯW*$��s�x�}�ĉ���;�9&u d&34SY�	p�T�~�Nl��a9�@�Y�1��m�Dn���S	��r�Uq#��˕b��J^��zOO;�������*�|�R��Bl�&DP�%5�V�����@��D��VD��W�I�A�?�<'\e+�ٙ(�gU~���̏{{�gX�(Pd�sg��=�*�a�*t�:����
r���eM|�,��p��ԫ�R˲Q�	�=M��%6�ƭ����7�]�E3a�<���'��&b�$S`%	B��QDeg@`�z���6j���J�^~r�d�M�,��[R���[��%F�A��FG���̷~��;�|ͫ^��UW ?��1/�J�Ç�>x�=�~��5#���*T��r	d�b�2�n��G7T��(�V�0����M/~�c��OL�����u�jsj|���_��?��W���{���_�����;L�b=#��yJdi�\�y�����W��bѹ���ן?5��'Rz�S���l����5~���Q����!��N�ض�%�ܘN��q�=�ٿ
�~�ݧ�3t�B��E\���"�q��x.��7��W���ѱ��w�=td�v@x���V��܅��5Qt8��2�,1�tؘ���}���ɓ�T(O�^��(@�+�?��4rN[�D�j��e覛�O3x��(o�qP�u�V)�tu�����y�������h�^/9>r�C�/ٲ�dz���NH��5�d&��b(&��j�0a\8g��H�'�i��O:|H»�0��Ĵ`4�VF��"�9��h���>�^�=G�D@�Ȏ�E��H�غ�iJ�EH3����Q��G$@�wt�����$D���S�^�% �!V,%�>�B���kv!���K�A6a|B��t�$�썠1�j���!sL�1K��=��?����&'��z�&���[^2�f�Q7�E\c�Pʨ�Zd[<���@iy����ٳ�GQ,�E�K8A_���O.���P"K$�Y��Z�MM�=���C=W�`b����O=����^��/[M;0�dR�>5��΃O>yrl��R�{ggWU&���k�ړTv		;T@�{Z\P�]��U��E�ݵ�G��N�8��3JϨ0�OE!�K��=�Jj_޾�o��9�U�����&�6]'�����s���9�����u�0�#�K�#��� M.�b6`bj�;p���`������    IDAT�BP��l9j�����e67�C�>���ݒ�GҐy����� �j!@WDK��TADlM'r���d3$�1�͉�oQ���"���
��[��� t���_��ug��������޷O�.�[e���&��XHۄBX�� ��_����n",�c�o;4H����]V'�
��0�5���q(9D2����x,G����dRط��X͘�|���\���Ղ"5W�΅KīA�$��t�uX&�U�Yb��7m� ?Ab%���">�QBD�ҕ��	�K�'���|��?�y0G'pr,�v�ݼ�F
�5�����cӦ�3����$v,1B���<tdׁC;���� �9�YD�)я�qT��h��Zl���C�����5�#� 1i� ��P$�P ��SẠ�1$5$*ƲN��q��sEߣ�AAK�]c��N8<,K��6 ?�
�.��ZP��N�m�A]�ʎ�.�����R��t�`��������vݵ�6*�!�*Ş��|xK_�R�0�=���X��+;��@A^2l��-p�C��GF{z;A��D�9�38��R�d%�H�TI%� ��+��+���
���25Ac]m�p���=��_�Nf(B\�k>$�ڌ��D㩸$.4T�89�;ԯ^�d,��*,A������v�c ����6]����X��!I��x���[�Z�ȋ0�56��64��H����8[��i�$S1($�E ��)��e�FR{��'E�s|r��=6{�dJ�X�T�ڽ�#�^9��"z`K���$_�ȁ��FF��񬷔��Æ�|Nҟեô]=±:9:e2g�D�I�q|��'�6�@�9��cՊشʰ1�T��󺖙^A�KQ�i�Q��qƷK 8��8hxh4�E�yY������+5SgגTj����O�8�,�R�Na��� h^���0�M��KN?�LP'�	�+쥔 ��DMd'7��XVN��!�B��=f�QL���V/�H�[�#���¶�"P��o!}$��{XD�$�;kަ%h�Z^������+��=P�����[^?Y�3C$P��Kf/i�dQ��>_��ܵ{2�#^-��Zyۧn}����8 >�h���w�z�Z��X�-��-q�ax�b�p�e/�t�����ݻ�B�B�c�!�D�5�Y���z�s�Ĺb�9E%56�GF
�A�Tt�~xG�j�g�RK.�)�7.�eռ�����C�R�K�I��g%o����P\a�1����d�8�V�d���7�X)+cn�f��nbn�c�`��kN��@:H���#3�Nl\�/!�"�'��6�*a�hvKH�̙��X���f�u�D��ʆ>��~�+>�dDC���)2��ي/qQ,�JP��b&�e��8��o.8k�[6<�hlh�H�¸9���X����Ӷs|���H�f��+�c	�"����z���N� #��i=�v��@U��~���&W(%��ye��)pf�$Ǚ���L3�b�h��\N��=.����S��_p1K�m#�̌�`"�
�'V:�\�|%�$��qf;�qLv�f,*�� p�E�I�'@���2ۖ������S�L*p������*UB��J�X���j�=����^p��
�����IZ�x��V�)��Y��\a��ႏ`�XD�\ SHdx{�`=2:59�=�4^p��9{"d�L��m�Tk�W��B�C�9� �_��&b��*�]�.��Ӕ��K�g�����Y���Ofk�tm���+�8��>زTAr�d$�7�@Х9����Q'|��"a�D_'�
�C�I�r
�nN�:���h�fV9���SK�Y���c����DBr�r�E��KL��L�d �J�!�I�� R%(%�ꀏt�	�ݣ��J�(�uv���E�!���dpAd�\0��*���1�3�h,�a����7pl'F��ߔ0�`nUk9�H�j�p�T�~�r6��NM��G���._�K��.w<I@ "2 �Ӹ���ь�5�N��D,�t$b ��E����	L����p"��D�YM�՞K��N��A��B.���	���]ٜ5Ԟƨ���a��4�=PPCĎE�^'e�^[C��!��?���+������A��ae�㋙a�� �"�?�Q8�'h9�#�MI�
�l���C��V[�c�f'�l�3�^�RQ�H��E��j���Nn}��w�h�I�p�ut|��r�b;m��R��2P�evK�J�
Ҽ� �Q�����^�*@�eu�E��+�j�P�#/����ʖ���˖-�&��Z�\��ػ��u�N �G��+-�+�T�L��q�;w��gdxlH�O%f����Rrc�N7�-MV�� WU�E�7�(��uY>��^Q��[C���$<��+{��CԪ�6$&�x�C���W�z��:�<2�XҸ\�ǎ�����IQ�3�Ej,xS���q"B�=��Y6�X���j9�W㉂��T�"��;���������M>�������|=˒#޼z͚����bmq{����+V,��:v�O�9t`/���곷�4
�4�5A��>^4 �O_RS��pY��i,=!V�� ����c�)�=��;n��T&��oUw�l�*�&!0 �(l1ڐeV�){'����F�d#ڵ��ѱ�뮻�#OED��wg2Q���|�T*ςI��aX�ׇ�A�/�M���xl"z*.�S�8i��31�L
	�#N��K��ډ��bX�K�bn_O[��U��a�e��0��C���r,C�zQ��z���ԩѥ�"�Υ���X�hl�1�/V�Yh�^L�!E18�]M_�C�u'H�H ���7W*�Z��r��-���������BVf�&�q����p��Y�NFF`(���~��M�uLND��1�&F�k�P.�Bs��梖���]� T�Jo� H��h�l.~[�<G��h��w;ۣc*c���T#XZJ�Q�	�F�B�
n��q"'���*�N��r��ys��X�q"�,_��-�݀!���D���N ǵ,/�T4�Ȗ9�J��y��|��^N�$�J���숈��F[sӜ4�eUt��uxyN���/��?�k��x,��{��u
 G)���A��E��"���Ʌ�"Q��v��� ;���'zh���ç��T����%�K~��TkΑ����뢱DAb	��+Mt'����]���R.����N;�P�v���[�{����.������Ԕ4��eqxZ�/������[^��O΃�=sӺ�����8b�"� _0r
]�� t�rt��ꗾ��1I	����l ,,ٽk�L(��a�c�� ~g�.}>��%]GF�n&����	_��7�Ld���֬>���Xv�l���N�����k�[��4��1009&ǧ\��h"���0xs�*T�4�G�b�ԪQ�����P�-����eua�$�k3�1K�C�L��P��0:�g�R���!�2�10�7Z�I��k2��ߗ^�i���P~; �C;������/���s��
�� �hX>x&� ���v�F,S���� s�ZE�"G�d�=�/N�!��>1�<t`����}��W%��X�pH6q��ܺ�"�j�EFKٝN�8 SnA	E(�D(��T��O�]K��=+��s��a�&����G�$bj��ٟL��EzӪ4�����|Z=�r���	Ѣ.��缑?sn-ti�~T�s�`PF󞟾�oOb����X$s��u�1N
�kR=?5GC ��y�:��"�`��;t%C����4������۾���]����p�wI�[w|y���z���|��=)B��ln�����M���d	fsP����]�(�����X��.u!:|���2C�6'2`R� �> ��u��A?�r�R��V0��(d4�������ΐ*�[�	���%������ ���9� S��z��r����<Jf}��t-��	�-=4�y䡇��W�fr-FJ�I�|{�ȓOnɦ'^޳c��H^��#���J-�F�j���M�����:C(L_|q:;a�b�w��ɩ����5��p�On} �k�j�R�LC��� �Q!����|����/��P�1xt���z���OQ��XN����W�hQ�]�d�י矉!iևG'�>���C�v+�1�*hZ����`�����"g�K��N+�c�H,o��iko#�>>CC�x�AM29�P_ȇ�f=��b�X�1у�6i�IN!�ۅ�\�����W*�=�If<A�D �=T%j��O�0���.�����N�Q_��$���7�%mw�9I>��>�q�!�&15!�A]f��~���5�>�]���i�~e��;Mc򕂓H�����J&���޽��d��zĚٻ��B�S��rVa�Oɑ�m(5y54%ݔ��T�d!^�_�A)�G�=���;���>?�*������#�/��'���V�_mV1� S,T��-�ZVE�O #'RGa_]��
�"�B!�@�]�LX�V��3��������m��N΂�h$�M�MƞkL4
�N�O���
*������jF���"�A�KA��2�-t.~B��e�E��yqY�T��Y��������hx��l$:�I���S�O~��w�E��b^e�h���,��HA�#C��o�L��2��L��KG�^.���"�,���~���SM9 A	�mH2���/E�1w9�|��~���C�Tܿ�E~�(�,��9���s��Q��B+i���s·>�w���S���&w�܇�X��pD� j��D��f�/P:q9a����-1�?r8��O}b�s[-6�5��C=#�#��%���Y���B�VD]blL9p@1�LM�"@��j�YJ�^@T&�iZ�'>q��>�~d�8��l������D�� N���F���O�J8�q�"#�b5j{��6OɋU~n���7���!>抳<sHU�D��s����	Dg��CN��\�cT��IYy�ʏF�M(N�&��V.f�-�+����J-cs�t�!Z�*�+������X���F�6a�(��hם�[S������U��ί\yv��kS�{}��u�W�1��X����P�;ӝw|�ɧ��r�=��p�''���i�1�=���&Y~����t�Bl�E�O� ���n&���x�(!�8��ʡ�T�v7b�\)�N�=���\�W򧄜½��ѳI�U�!�8�L�vCњq2�!g���V!ad"��x��X)�v	�.�GPd���m0���37�q�Ȁ����V���0KZ�4�8KT^�X�rPI����`]:��zȎT`z�fAĆt�Z3�q��P��l�o�Z�l�ˍ���G��T��*AY�E(oa�*4J�T���y�wO��;S���Z/���r�:��o���F�'�(pÊ�ᇟ0ۺ �6��1Ю1{��O�ջ騲F]2.Y��WI	�n,�x��� �zp�΃��sƜM4�><L�������tP&M)9�s8��]mł1/�����5�6�-@��� ���
��g�	E�S�D�"��6	�@W��H��d�!q+Ȱ���^�1L$#�|�D�N�ԛH�N��ޯ��?sT�^�rӬ��2Gxd6�P���\�W�šf8ӏ�:��W?}�s��4��x�}�v��(
�Y�W�6)=��r�2Z_<E�Y���ա^�l`�17�&ANV	O9�E_gGw"��7�jv����ů��.�=��1�Ϳr���ۈ�O(���%4	qo�ZBXW�����([��[jX�l�h]�E�Q8Q�Z.�&r���8|���`��Sig��/i)s�Jz]8�r!��N�Q��H"�}|���%6Ie!iq*cj�~?*P�U1��VȖi���(�D�}���-�Ã۶m߼�ʏ|�^��1�xe�02�B(ԅ��e	���'�'N»+��l�c���2h�tW�;��c�?{� ��G���Ϯ}�-�ъ I
@н� ��:�*nw�141:`�@�4�09{�n��z�5��}���p�2�����-����'�m��<�Q�Jh�5��e�5��)�RIb��"�x$j��A@�%���޶�)���L%�^p�������w��<��-��탉�D)������p�>���7���5�ox���868�fW�$����K�,G��d�>��]J=iE��b�"E'P�IU�;��*\=L�	���y`�Kze�"���f�����b/�����0Y�q]�����\��[�j���U����
ĈL6�����Q�{h-J\O�9GP˜+������ d5)����������b8�ᛙ#�]�g��:�Tc�W��	�R�o�#t C�%_͌��\�����ޱv�W�q3p �U8�&'����5�Z�3ڜAa�s, E�/��K0�^�
*��*����HS/��S%%os�ӹ,�Vu5S�͕$�- �=��^E~�����۪���N�cW�G��㓤(`��3�,�h��y�uA�����d��ٴ*O2̙L9��g�L��e�լ�)
t�)�R���fh6�ĺC#g��K����p�w���֭[W�}�e��r8�k��qǮ�-���BU�XS�����%���a�0�($n���W}^��#bժ���\����;x�ޗ�>���ή�k�$xE��,���R`�v������Q�t��k����Lg��U��&�Rd�볓xd&���2��"Rt���r�M8���合W�F�q"ܬ�-
*���0�GG�o� �%ӡ$bp6C�=P�J��3{S�qї��]q�E��ٻw���x6o�a�a	�Ld�\za���������)��4��c	IZ5E�X ���	��G�xbV"�b�[Ȗ?H��ő�\���@��i���@� xfGf ���d�w���P�i0�u��x&�Z�T��3��iac��y�*G�Ð���}D�6犾�����e�64l��R
X���v����HZ�ґ�SW�]� RS�/ŐIT=F����]��H�����j�E�c�=K���w��tZ޷z��C۷�E@��s��$[r*�T���)�+ tb���݁i�6hZ }��SM��򜖁��ˇ�f�6Kt F�˝�d>��e�A�c��d4
A�����ċlD�EY���͛�Y:�@���W/z��]��xBd6���~�g�={S�����_|�C9���T�jE{��;�Cp�L��ԡ o��0]��$z�|����a����'��&ӹ���ۻ��_�����'��@Bj���&�	hs���'B`%�U��A�b`����f;�l!	Y��H���tS}=i�+!�h�K,��=��
L}ح{��E�+@w@Z� �	�M���2aE�Q(V�$cg���]#�`2Q Q���Gc�c�M�75j��������d�����H8�w���S9��T���׏�<f�2?zQ��q���B԰M_8%'�JCpb@�/���Zk��`�њj����9G�|#�R(h!G��9"�� 4��D_�=���k�K�Y�d(]�]O2i�N��"A���l���@�bR03��A�Cz��\9!�nǹ睝N�v����?�8�dx2�i[��3c��d�M�b���uJQ�k>ȕWG���V�3�as������H~hH#'���tbxh2�#dB�J��1�KB�T(zz�.�2�lB�r.Sп�������!�j���8��9�����H�6�#�`���[��~���S��;�v��g��bE��'J[�yBqÆ�Id�b��/�dg"�i ��نS�� �K{ȹ��t;���؆�;Ñ�������#��庫�y��x�z��xT�V�P,vt��S�&@D�����ly�UWm&EZ.A�sh�$�M�"�iu�ޫ���v�>�%�]\�hB0�{��9�B�͝��&D�,�ؿ�
A���Ϫ� _P��    IDAT�>.��&�'�<"P�L����Y�	������]�$�))^��LkV�T� �"�C�%:�*��H�T��=6�[bq���8�=�]��_��~� �T��;̪p^b�	�ŷ+�ŧ.=�zd�e��9	��.��L^`Kt��f鋴HbK���Q�8B�ԯH<�F��}���\�R�k�7���8A�q�a:69Ft8'�9L^C����.q�969��b��gs�1�M�ۂĶ@zok@l�+(BMQ�g5����R�C}y�-�������X��$c��)!]�S#�xT�0y����b)�~F5�r<6AH%_�� &��ݐ+��q\���m�z�i�"?v\D����� ƄƎ�=����G��/������O�/�~�3��/ |��3��169I::a�UIXlrv���2�$�?�|�:��d�:w<����O\S��	�z�+�p/I)�.�@6]˓" ��u���hd�~h����n��oI�K/l���ڿ������)�ԍ�L���a���߾��ǟx�~��[w�x�p��Bߑ�L
'�1[�Ӌ�Y��Bz�LN�-#���Yі�p@�EzE��+��П�@5fR��p�y]��PQ����4#n+��R�b��"�8xldӞvӳB�Kj�g)�&x�,UXV�-Q܏�Ԝ���Ғ�t�^����;u�:*xAw�J3yF��B�*x��j拴�gM;�z��������!cD�#�Qm�()�X��c��v wH$���Y&�5.���5�1*ؼ���u�L (�ɘ
DS��A�@�������^]"?�T����n<�:�x��
�L��h�L��6�m1�b9��`�������^��u�@(�D���[qVJ��-S��1-�R�hU����=7����α�.��:|t����-���������
҂�-�RZ�PJ�y�:EB���s��W����d����%�iʜ������=��CG^�F�^��=,�b>��!m�1�)l�~xv	Rº�w����on������7� ���4Y�b��Z�x��$X���QU8���<*���HV�>LXĲ�Iё�<^k(�$��S\�t���Q2�}�4<n��+>olU�4��" ��Pp�-]m$x�}���#����[\^���ށ�a�xJ�K�Ӫ��#YC��(zJ��Y8��ꕼ�S֜:av6�]hkdw���:�eg�\&eAG����L��(S�)�#�fLL��Fw��?EG!O4jVmP��pX���.H��F�V<��!n�x�r8�����6v���_8Ϥr�j��p�qc��/da��'�yFB�4��o���*�i�ob�Uv�9W�T��
b`<pd|4<V��4�ں:6_|�ʕ+/<�\L���LE�߶��'�:x�H1=5����%�V����G!���
ހp0�M�d��2	ev�L�_�m�#��4�u�p *J�r ?�	�{����i �%�kӌq|���nk�D�&
��Nl*Iǂz^2����i,�!�-�A��1n�Ǌ�f���{�!��C���(���!�$L$��B$:���\��f�PFP�uQ��d���?�ܻ�0O��rz2h��R=)�Zw[=	GzĦ A1f�ٞy晏}��s2�8� BR�(A�5[���d13E�(�$D'��`bۑ�=���d�,e�mk�,[��y憾����x�I7� �-M�/H�2�2�B����lF�p�핎v')C�:�Rx����������_�ȼb��J�<�:6ݘ:�` ^���?���D��Q'� Ƞ1�h᫟��0��3�r����
Y�y���SX$�f��Wɦk�v����prl��%� wǅ����Cm��D���2>��W�y��G��)`;\V��O@g���r����wHO�O$fӽVo�3_N[n���A8l��&|��%\5g3�������\ұ���_�����eK;�l@~ܚ�=7]�w�}�x��'I���'����/w�TPE�%�@��~��ы@�AB�H��,S6�y��P�Q�Y��\*{�#<��\Y�����}:�)v�:��ߎ,�s�:��vYWy��t��g�\ޖ��r�(�1�d
y�Ŕ�fs�9��:�w��h�x�������g�;V�01v��jt�� 𛡊��A�0�]��bW���6�X����M���PL��*�SL**ʙ�L>�P���>yER��(u�~�d��ڹg��v��gs��.�t���-ED��Gx�K�P��g:0D$o���ddr"�
;<���c�b�4)[�~��_��M=��rCR�*�aD����ȴ�Z�;w�>��K���O>v��N4��x�h���ɩ|+1�ǞAYb΁3��?QbkN%��U�]�ƽ��e�� �dC��LO�(����n<q2?OtR@u�W�^C�v�T7�i |��"�5%�)DL��S�|�b�2r"�T<<96T+�^�9g���w����߰�' ��'�t�%Æ}k�����{x�M�O�V�׹<��B��S�T֧�ҵ�r��\l�/]R�;�҃���L&b������z׻����t֦�0�3KNp�F u��.~�&P�/��7��o{��8z�Њ5��e�Ϡ^'�ؐ�A�A�	U�g�JFh!5$(���D���qT�4s�Z!�&��!�3;>15::N/�n[�h�'p�-���h�&������|����z�U�j�hxll�X,E��r�F���H��:��s�K�sp4�|<��5xl"6Yz��������=55�KA�� @����Y��V��{� 2�@���;c�:@O�:+DO�p�,u�8h5��sDV X!�m�l�c1��f��"��'p��j4T{���8�#�Q��ȗ1�~lt�)���hJ�419��n��L�HEr�=�A+,<\�'2��f������Q�;O芜����hY
��
��,�Al�>A�@���_}1+0p~�s��8������0��P����2ݹWO�wZ�*[�Qɤ�m�e�4�U�g�R�ɆuJa���G*��!t��_(��U����ћ?p�y���|���XoH�ogu����/:���>����}���p��o� �#�]�:d����xLR�_�|2�����O1;+%ɘ��+�I�&��N����9+y�jS؁��O�Ǐ����n�����_o64]|Lի �Vû���Z���-�O��{W�Z�˖ʲ��{�a"��WQ8&��P����O4I0�@FX p��R%BX�B͑-�<�n�0&����G�ۢ�!Z�T6�,��.�yo�����b��.Z��<�X�b/x�)k_wg��G�V6�qŦ&A�6�����K�|('IV��y J�Zb�/�� 24����db�B,��g�,N�Bd+��n���	����/�cf󀌺��	&DTlN�:v��h,c�,���J􈘥�'��T���Il^�`R`H�U)c�ML(���t��.���#���*��X�V�&�=�%����0Ca��JB�*s�B�\�N�ˉ+��"d�+�LnK����{�t'�c��5RYQ�'�T��Si��{!b Z�6�u��i-�Z*���s%�:ZH�|N����{�kyBO�˻~}��������u��	�f�7'������.i,�rG��h�.�-^*N^��k��7���4��U3w�V��e�V(Q_�����ט��o}��{�"�=�$���Z��ƉZ�M�}�`<���J�v��R���R����Z����ۊ)/d ƒ=]��X��< �ht�z��対�oY����OeT[G�u�΅�믿k��|�K�y���5�i�X:���˶�D�έc�;Ph���!aʕ8I�;F�U��#U.]�W|�DE�by��}�������@-��NMaC2�͛�dr�b��ALܹd>��X������;�S�o�@AN�=�H��j�X/޼�7_���~��{����>V�vQ�-zĀK�R�|`1���ܓF���#-_��#��Xsid=�7]uݭ��t�<zt�ᇶl��"���Iw���ѐ³���Zz`p��t-v�=K�����M�W\C� �$\?�����D�Hc�G��.���N����&.�TH3�9����F����%�gWe^"�����ר}��5&��N<r�X|cc��1��~��_��gV��a"���2��4��e���}�i��K�?��)�8�d�&Գ���,��e]�S
�d�,�)ȭӄ�^!�U�$	}1�A�I�Z%�o�喛;�d%0����L��i���Xg�����iˣO�'�!���Z�2(�A���WU����)(Ds=MW�"��B�N�3A��\#E�_�B�8�8&erS5b����@d�b�H��I�-�"�k֢�CqLN�R���8�q@�ΣF�C�W����'&E;nB6i *L.#'T��Gd�e�K�o����_������O��:<hN@ք%#��!���Iy�+-Q��Ax1io��J�z-��2�\�b����8�0l�ց^�(�5�dtI�u�MC���x2�
����ۭ���'Kd�$"�K��Nx����I�^�E�ב�U\�R��G�]�#DS46�.�>�����1��d������R�b�� st�sļƄD2��t��?���+7bY�����.ɦ�����/x���n$|�\r΍�zǶ�^�����'�}�L4�,N�?B+�C�4�K֥�qS���5�LV(1�h�5��G'FO[���_�B�{u�Gc&��:��6k��޼ȥ���f��׿�u���w|�S���X��4��!lB3e偲�"Jo*,{!������L��E�K��Ų����m� ��
Idն��-���@�L�)�M��pZgOw2���[�uǆL]�b2�tm�D���x�6�1����l��`9�[�	x+���[���*f�\=U�D��������ߟv�{^���/�d�O�ޘ��>�)�B
����V�6:�{ �f��v)P�à�\1�����n�����򽤵-O�FZ�ġ�ϟ�6E�
�Tܜ􃎋��f$��K;�����>��H�2bb ~e.
��K�J�)�[j5��Nʤ�S��4�*fA�/sR�p��ԓ�G�I�P7hQ����nipI���
���Zr��qth�\L������z�E��u,���8C�S�7��x��t�;H�}���O��*�Lx���PuMC���Х�����,ZP ��<ǎ�-�$�|*�^w��gt*4!��iw��iͬ�����R��=���&ҥ��'�\���\R��H����$��,���H�~���x���0�P�,E��b�nL��PE�R��b���.Z��ƶ�qX��+��,����p/EE� gm"��n�j��T�P$�<���7v�N�����l���������T6*9�6N��GR?�����Ik3�9�1T��������,L< �?�|L@xTUl'P�`���V��Ҷ}��D�]mm��A.nq���$-���튎���!�+�u���|�?�������ϔDQ��c�d6Y��G^Lp薍�����B�T1V�R�B������d����l�$�L���>���'�����e�DF��
]���;��z�W���� s
�8.�D�1[�鄠�?��7_y�f���DX�� fm���[XP~�7O��O��ޭ�m��/~#9�02Th��+�l�6LW�Х"�}��Lcy�;���$"$����������{��4�%fS�Y2I����޹�	N���|�J=��7����?0��/$h'[��^��k��9���O �z��$KO6�$ʙ�_�^t��^���H��T}~��/~�˗_v��o=r`���0���#3�=U#12,�]��է�c��߽����'�5l6K�d��P��׼�NP똣J�p� ߬U�����!�ǞI� ~������D�N,?jB���^�Qf���#�ua�\���md�X�D���.D]�6�Aj�����z�jl��m�����淾�"?��СC�>X�k)H�Z�	�m�i����H4l�%W�3�3M>�U��	���B`l"\�Xܾv�x�pQ?3�{xP,���35xfU�{|�%��S���3@�f�fR�����EQ9뜍�l>�J���*I0(�]E}o�(�w||t��^�|�Ⱋ/���{�c���Ǳ���x�)��Es�X�j��"�N��x=<�Zp���ȹ�	M�}Jj2���x��_����>��#)��.���(0u&K`�Ob{C~11�S�w�}���|�o�K�{������t ^Cf��O���!G�����9����\���ѩ�=zt��ͷo�)lH!�5�ۓ�٢�]�g���{i�5� �+���򦚷R�[���ɟ�,�Et3Y� %*��0I'�/�����v�ۏuwg'�qV��]ط7��e+�^H���<�%"��Or�H�lo.� 6�Dc�'n��p�f�$8�wG�Q"S�a��*]�x�Y�+��.��+�NMfv�E�c4��!�]&��D�o2jR�4$��`ו�D�T���� ��$�ۻ���!d!Ymm$W	����E�@e�\���k
D��[��9�ғ+W�}�������&$I]�:&��f����bJCZr���"\!�ʫ.;��s_xq<61NV?�a�qb�2�gף����.z�jM]��(���VK~21�y��^vQ2�J�k�5�+�H�+!o7+�\��Y�7���@�xH/�[r�-���G���6'i3p�t��B�0���۠Tg���o4CR����8hb�7�M��\�����=���b�O#a ~�� �Pv4���u�;x�U�1�!@p�݉T�����^�ކx���.O�)iud�%� &��4AI��2�%�P�/�◢�?�A���LV��tx=~�d��^�g�"����E ��,��yM}ǚ�:2�{!�aX	$�����?�F�I���i<���D. �ta�u�:,��py�#c�l�����?��t����U�p�
}�|�$)=����	u�Հ����~����� +�d�F��ؒ�ҥN�p;E8��ȧ,�iX}��n���k	,��ǓNL�7\�aݻozG[�<(�8�阉� ���,�l��ބ[�\�ho���̺uK���w:vw2�d��t�cިР��̮�:g�K�H ���R
E���[��:����\v����(�W�@��
Ñ}f�μ���DC�����i^}�/������q����xo8c��>Y)-�4�?���b$s���g��dxh�;�{�����e��|��]Sca����̒�">�@��M�J3ɂ�y<��H�L�T]8�Q�ذ~���L��Á�y����~���6�`��|�Ɨ�a�X��E���C��T�$j�;�]�;�&��V�XF��Q��@�@|r���lU�K�U�ȃ�P�&7�D�,v~���ۻ<5<m��(���WS�@'�i�ޏ�q9�A�,���wzLq[p5}����ԅt=�t����t{���n�_s��^��	b�J��Y��������@�h�]����U������+����5y�����nXD�b1�ֹۡ0j~?��"q=fq:�O�֘-kQ1�I�� b)�+>>xUD�?�o�s�l%@ъe˧����Lgg'������lwI85�'���ѐ�F��H'���+ɻ�g5�#�/H�U�5ӌ���s�T¥`�o���ۃ�`���*�q
���j��d}9�y�MW�OD��mp'�:y�ؾ}Xi�e}�Ug�]�?hmO�;�/(� ��'�OE0n��:!�lGe�,���I���U�ʪ����ʟ����r�zj��?:0p��9��n��	vN�W�T�G���`O�t�@6"^[�_��_���<rb�@܉���%�X��DAޫ�(  UIDATfB��u�^� 1n���.
�	ޢj�����eH?%C���l��z/T�~�>���J{���6�o�WG�C�4T�w��Z�x��
�D"�C��R�*��	��JY��"�?��7������)�� ����׷����!����J�Z:S�f;�mf�.3)!�8Uhެ���A�d�T��q�Bp��u&����Sk�Ѻ�ͯ��壼�$�Hg���e'Jc��b���2�)&��b�`���R=�0��O�P���D*��F�v�J/� 8�E~<J%~���: ;+L-T<�Saթ���@�A�+�"Og���r"[�]B�zC&k�D{^> -n�� � �(�]!�����QЕ�W'e����h�b�u��~��N��^���]9�3:��P��b$W���CHb�X�5O8A��E�\}5�e�G��R�v)��B��r��Be`sJ%(� �O
eW��D9]"Pw��'��2��(M��K���U@0��PA0�`(���!���+Yͪ��3i���,Ī��V<�L@`�Bl"?4�r(T�}��pjF��W�=]55�,i������s u�wV0r@�Z%L^,�}�0_v���B�ܦ��i3=�� D��f��!0#�4XRB�@��"&_�e��$��jp4�E^�S`Xj���߽����x{�D�Z��E�W��ئv��Ƙt��`]C��!q���4�>~a�F�bE}��DV�屛������K���vyH��Td
�� J}*����]�b�ф}��BY�T�
5�dg�S��N|�#5(t�+ �9ʼ�t���w��1���3��tiƕ���_���A�I���	;3G]�!���K)�p�9Gx�E��鲚�
Ъ&�ƋD�X�g��q���k�#�07�-N�MC�|[��g��l��kl×���x���` w`��:\�iD�ŔLa�'�Ik��o�y�q6�.�B�����U�xLv���x�P	���)C.344��Lǝ�
��?Ռ�نLj��o�(Y�Α���g�B��&�z��Qm�S��
��&@�Ta
�����pV�����a���5�p��\@�UX0�ݝ)��	�tNQ3�5p�^��b�riap$o���X���E�@O�B ouy��ږV+���Q��KxPᶥp�yH��bޮ�-��r�
�TG�V���/r�X#���O��+���S��Js	Zf�p�+�o��>����f�lݪ:��7T��2E�!�f7 sI��%J�Ю�10h��tW֯�A���#]IB�cbQPo���ƀ4i^�ݚ;�k�dou;�Q�� +�{7���լ�S=�g�~
��~�D��4�L=)[2���(�>���iUf�KM��Y�����p�����;c��B�s�Xcu�
�%FՂ�Xs��?��-?
�8qy��X�w�{j��k,���*j��'�fn��=W`jVɂ�}�(jYwvv����H2���h,�R>�M.���4��D,Ո���c$b $w�+��Db�N!�7,�<��~ qC�fCli13������*��TC�����)y02��G���E�3�/�h�	�.�I�Q���ɴ���ܽУ�E�'X�~ƩP�
��/ {uEa:yM�P�m�XDLLjQa�&ʆ�%5>�-5F�G�C��T�w�>*��qW��P%j;���� N�� T���@����_?`Լp��y����'�V2!��Q����A���N����%��L`�܁c���۩�	ޑ�ı���+����A�X��K�4F�	�.+b�?���r%���7�a�$��Jn�ĺe
5H+��L�t�<�=)��d����}�P?rP'6�CBn���NY�󕙗ʽ���-L �'�t�<n��>� k�h��@bQ$Å\䆒�PXTe�'�g-��D%8�r��9��tX�6I���WSv�lrT�A��0�BB�	�����Ŏ�"X��>��S��坼D�[���������T;�`˦�"��p��e�H8Q�:� ���ߎ�f�`��E�?z!j+�S�x��XW�%Eڃ�̾��~�=ĂE)&����BB*)�j�L��y�Ho<����� B+�ǉ7�s�f?|��[w^|�YӚ�z��3C�w8�����=��0�Z~���'''�^�L�z�D���&��Ȇ�+3�u�r�CF�+�Ɔ�9�ȦW�^M���ѡ�Z��d`˖-N���V/9������A~�7W-P�����v@K�C�N	8+�w� �	��J��f��|�2	O=�>a� ��9!zb��I��r���LD�H+L6��H1�q٩� L�D�Q�9.,25��i(y�)K�`��� �t,q�������kUk4��x]�����0�:��NDvR%���c��/�#�=�F-D�r??
�&eaG�/�G����S?^�`�������t�eW6.���H� /I��ޤf!�j"x��Q�� |`)6h�2S�&�딣��h�T���!�g��<�u,~�V!�����l�v�ޝ�~��[����߼ɪ���pM@�^�X�XmV��D��{�TB������/[���ͻr�r96-��:�}����T^h^��֏�����}���X�����l��Ԁ���h��F�n����o\w�a{ل��%�!KH�²W���HR���&��X2x����eN��������n��41kTv(ʡ��&qd��7�D��B�T��|�$���a��QA��!�H3]0�-{Dm��բ�sJ�y�/�t�Ey�t�)��O�B�+�ݏ�c>��㋢T9�����D%Q�,g���3F��f�rj��UOg"0�74�S�y�, �3U6��J<���G!\	�
�0|�vcU�<��|=f��NL�O|~�N^���JU/=jB�6�\�`��z`����N��#h	aĒ.�2w|��������#$QD�F�4\zx��0Boز)��]�"QJ��#� z��CkR63���W��Lr"Zk�3����]������{�&����0	%�j�I�	�4
������zCww7�v۶m0�/�x�R-t�vW
�����<��s�{ύ~����Sctr��g�`Hj*�c��� T��D�e����j�J��J�����~����A��c ������`Y��
��s�C�sE�#����h��W���j����	��V��������?���S����ϩ~�b�'�W��	�]�X�<(�̯�Ѝo{[g������{�h?�)����a0�\0v�׀�	ڱ����zܑh,uu�=:v�O~�|�qQqL���	\{�5�6mB{Γ�͎��3�_����Gs���x��}��XԹj�꾥+w��i��	:����s���_�"5m���6p)�a[(l)��DQ��,�b��tZ�Rv����|?<�������ا�M������S�%�	EcP�G��k�7_W�!J��8·�$�o�7�̖휯��}Y<?	��'��ٸX۩� ���$��3����@%[}�g��c�����{즑��+VA�v����VP��0�A*n�ҁ돕Ԅ��/ʻ��-?��}xQ�v���7c��K7_q���T*�kH��fP�h�򗿬O9b�I���f5�]����?\2:��v/��=t���݄ҊL�ٳ���֯w��xH������@�d�f���R!��0j����ٵ������l1�=���Q��/�DW��W#H��@�D�|�YG�e֕��XZ�����Ť^�-� ��κ����!|�u��9=�i��.^��!0?��:G���D��f2�YQG�m�t"~��A0�9g���ȑ����Q�e�b�#be�����6��������%����[}���Vn�Y}�B��z���ٕ+�@�
�6��Bz�i$G0g���E�#�����^t�E�^{�ϼ46��0>Qok�^�fM��ɉ�>��T>��[?��� �5�f�E�)"Ot%b�"�8쎟��;���۞}�@�l�/��!Lf�;#u����,��j�B���ڲ�w˛�H�Z���z��:�lt�m�_�ϿT��k�| ��j�|�Y���A��:���r6�A��pzq醑M�&���������|EHx�BI+�,�9�y�X�`mc7%쎝�����w���w�>���y��%֮]��oX���b��vA��X�0�3�%&P	;fT�Z�ۋr��CGʅ*&�$��ebb�R&a_��m����r{gO߲eE����i&�D�1��J����<�����<�o|g��'J����Q!��hj1(�]e�����U0憐�~��"i�qG�k��t�G��T�d�:jkȓ�Γ�ٓV�Ƀ��i�[{^{#��٣��^����Jv�j&ѝ�H��Bv玗v��ۻl)���B���P�p31wT�-�$�:)L{|����������b�G�ƴ����U�7���o��J�ۙ˦��	B�)�M[�	,�^�	�D�l�j��ܰ���ǻ�i��Q����=MO�'N+A��gȥ�n���\��[?���τ`-�26���q������������~@��l*�YF��d"v���Ca�,����i	�-�|R� ihU��;r�Ct�n��Gq�iU�|�9��'z�|������_��ꗷ�����U]����ڿx]C��`�Z��"�v�D#�����y���A�ːO����]���~a�ʕ>)bĄ+B��`03:�ٽ����|�@,D��3�~ƙgTJ�}��R����D\�`�Z*#�$���+.B��Xa���y3�p%�ց��m��#��X�����F�����<�0����`�m`���]���R����ɉ�;�q�Ҟn�?].�aw�Џ��yj��?[,XX�=��enw����T
�H��G6��=!ޑ�[���V�\!T�1s�2������W��"�����5�J�'p~\��%p��h�|�:��	�G����s��X��,\}�LR�r�J�X�-��wvt�/^���ccGGA�%�#�~j`��|��V���N��8�S�b��wo��忂 �@�ښ�ַby$<f0/��/���	���vl�*����+U�%�*
�4��	�	�x��_�z���^�P��@��������fK�"�Ap,q~KFbVb������	]��p�}� A.P�H8p"��.q��%1�l�p�ly�<�-��BMj��a�N�lh����[�g�����[ÿ�D]|�"� @$���r�Q18�G��	��ų�\&C Hu؆�� eW�P�Â���)�=]��rn|�h���V�[O|�/�>U�$^��T�ꠓ54P��	��.�u����}?���綃��%���T<�s؉���e�����:�(cP��!zI<kUR�bs���C�M�}�*�w�H���Y�=�>�c�N�)��Q�]�)9���oUN���jY����P!Ц@\�w�:\��P¹9юH�YBǦ
:rb�h�b<$~՘��]n��.y���Ԏ][/�x��?���������ܬ���$5�	Ҡp�"�43N�hRT�6Te+V.�hC8>�:�T4f�a#a�m��0�m7:�!�٣B^w��GK��O�V	��wy
�JEV�P=q�m&�:���bL�܊�s��o3'�ʪd��k��>�G��4���o���X��+A`��[��U*И,�ºB^0�rXg�Z��0Y�Q��6����>q�ݩX��5�X�^3z�����/P�B��T�@�%f�V����?̃.u��t:��3Oo۶}ph4I��u8��$�9$���&W�+���E,6h+,.��$�y��G.�pK���ICD����ĺ�TZ��F��{7�䅧���jY�|����ŋ�X�@Kh|���qQ�2�fK�
�<���$u�����?�j���B�R-���`ghÆӗ�Xr��uW^��3֟&v�}ָ��6M]��"65QcٹH3WL�V����خ|���x<:���a����Bn\�n�b%��%�%-j1�%2��9���4�u�UDl�ͤq@|	�|JKsOŋ�cU����\���ih��q 0%�����錔�\(�Є���&�=F�Z̏Џ�m.��5�&S��}�[��jt�\+Nu'�&�',<E�C-ī__�9�����C�r�fA��uМiblrﾗ!�K����Q�x�Pʗ%ܕL3�#���A���z���#=�*~�Eq��qc�u��U��Ve~jN��:٥xP�*�Qǭ�]�����o�J ؆zG�)��A^�k5�$��o�"��n&��P� P~��R�d}�Ҟ��$%�Ц37�Ͳ�<�B:t�TR�.g�K5.�&�l�X5��务��R&ޫ�|u�Ŧx	�*�2��Ġ�&F��C�����hD�VI���P3+�j ���!��E��j)��`:�f�#��@�I&�$�
�>�b�(9�ȳc�J>r9p�A�s��Wt9ݎ�z�;3��	�QǕTG�x6���B�4�BŖE�M>nb�	9���I�][�P���R.�z+B�R�bY��"!0/��)�*�.��ʭR!�^�"d��@T$��*6G�29V�9ېI�w�4��\9畠�E��8�,^X��"!�����K�X��"!0�Et9�ųE,B`� �Et�
�Y�i�X����,�!��E��?)H��=�O6    IEND�B`�PK   }Q�T��K� 	� /   images/cd1eebff-8d4c-4172-8358-6f93b12ef793.png V@���PNG

   IHDR  }  �   ���    IDATx��ߏ$�u&��s̬���_"��hDZn��� �o۲��4���/k���a�w~�_�I�a�G?�����&�ZY��"���RI\��a�L�Ȫʌ������U]]���=�3��}+3�Fܸy���q	l��l�����k�?,N;�|��8�l����R�:}쾺w���=Q��O�A+�{�p��ݍ������W�컗o���4�A���Ʊ66VE	3�3�1 ��L���|bwG�� ����E�Mk��`�c�T�fK�<k;���. ��p�<!�ݱ~3M��5�����6 $�� �Il-1��h4�a7��.��$��)�ԕ $����9A�:0� ���Ա�x�֭��#ߍ6X���`�VA�e\�v:���W��l����O��TCn��>�2r�������yf�/�i绺�G7n�:pف7�x��4�8����W��*� p㪝<���ת[��������1p]q�j��]����󋴽���X^G�S�G]�X�}wkw�
9�nW��n�k�/ �_�s��?����l��2� |0����h~{��v�Wf_��ӿtܸj��օ�D��Cuk���a�l�����f\���X�{�u��?�[;��/L;���_����z5`�Ez�ƴh���K�H'wk�����bq� �`w¹=��k���=%M-����|��&�k׭#b�iD `㎪v� x4�̈��e]s"	�睙���6hѨb֜Ț�4' m���d�*�Â�ĬaȊ(pqA�HJ*Mt�5���B�f��^�֑��X�Ξ�� �)�8�bĉ��OeѶ����,���[7o���y6���!}l��5��=�ғ�a�m�}���)��bw������-(�)]�-�i�`5O��#	�[�)�w R{��;"4<� �6Y�������wp/D ��˽�ד�t��v�Ȓ�R� f��(��Y\�JnJ�.@�EʒR�q��C �� �$Χ��� ���vN��Q2�7L�0ClG6�����	�g��{��>_Mp�s���1kZ����m�J��I���%�� P�HM�XP��5�&��BV�e���u�6k8f�ց_�T�u6��*�͕@]��
��4Kpk2@L�LFU��Ɠ����Z�"8 t�� ��YNۉ���'GSG�G�=O4����f��� ���i&sj<�mQ�q�g"��a�� i!\+tЃ��`�Ľ�`����j�W�ա�\ p6�yE(*1��2���0	@Y�j�q��gU<;H��nr �܌HX��p
�.��s���$vD�E���;XjZ���L��Kp�2A��T�X$����@�DN�Ⱦ �]u�ZR��f֌����o/��ݽ���p����|�!}l�cUm:������y�"���M�tA�BKVg �v��dm�Q�	 (Ufi�j$k��y���q�j�$!x�����.$�<�@��N��I�R�Y���C�:��Db����8J�kEu��"ޒ�*�N
��)~��-u0��F�+}. ��%q#� A
 -w�<">`UE�zb�j0��J �K�	�]�,��m� 0� ���8����$1֛�L#�*y)��Lr
�6��+ `/����� �������o3g*���K��4j���fdB,p1#6@�0Aۗ�3y&
�uq3�A������ȉ��!3w�35�fX�laf�1�HJ�89( D�D,�Np0*7�	�
^8�1S�1�_��Զ`6��#0܍�����O;�����[�Z(�`"8;� b��#r L��;�`�`q5��s7V�����sbe��`'r�	�N쀁�H]�D��0�3�3��RZ�؅@D�09��	�n��@p����F7��0� ܏���Cs��2��R7���_Q������_�o�����gkU�6xHlH��k�P������u\[�e�n ��#��l6��t��z��~�����eH���l|)H��/��t���\�[��Vs�q��W��v߸���׿Y���y��W�~�P����E1{e6��f^U��������鬻��� ���Oo������ʕo����On�� ���6�{�h�s�;�=':�;0 i�"�Q�u��ig�Uv�ˣ<ˉC�jO��խ�LRp���dZ��!�LZn�"�V)զd1RmYTr�,�� b䦤��X3s��������,,Ɉ �F�E�č��؜� 5�T�M��Ɉ؉p7B�.�Q`!� pa 7�Hԩ� R����ȸa�ƍ����Bd��I 8ca�#n��HU�*�km��NRiCw(��``("mXi˴���fi�Nn��d�7�12KHn�q<y[�@��n�R�9�<.�.�Z���ͣ�	1س�XXA�P��!����ȁTc�P@ b1��"Av�����Y�FB!!�`���6S7 �X21��3`�&8���� �r�@@V%*���ЇBDH�F �b�;�PJ��>��/ڗ��9/��{� ��X���D������%]~��%���BVEd9��&�����Y�DC@D`n���B������!�CX��>�Q����]��n�q@���~��27�aC��U\�����/�'��ݳ�싴XܦU_���6��>���C�����Rj�mƥb� �[e��>���{����lF7o~K�\�'r�������7?� ��Po �}���-��Ɏ5{����3�9�:z߫��l?���7��x�Σm ���6 pIw����kw�_�A�\�Ej_ݧ����+W~"7_�m�߄��7��ۣ���������ݶ�"\
5�٪�ȉ�N�|���G�Ż���&�CUo�t2��UK<χbR�w�I�B��#
 �/Q��(��S�J;��[ud ����/0Y�^Ea ��H͹jY�MI` �$�Y���)1��D�b�\A��8���ڲ����K��Y���q���q��Dn��T	lDfS׼��;3�AA� 2搌� �n@�n�pb���s�ى�����48,�A�M܉��9iMd�
n��V�1p�C�e^'"q��9P��R?/ܼb��j$��H8�~:P���{����rm� ة�O�;ء�B�@M���RO&�0d�I�	 ���ݝ�(lD���{S�9 �Q육؁�2�A��L`�
��s ��[���v���,�O�L0U���
���0@������(�
f'߫����0QO��i#��`�c� 1AXp8?@�����f�5"Z!�=��^i#�e�$h��| g�*��,�\U%x6dS1BX`pXV�	n��@� f�!<��렙A!�0xT��9�Ӻ��o�U���|�'����_�c�΁�&黶�\�t/��~�3����+s���6�?���72��?`�8ׯ��.��w��]��b ��4dO�J�/K�����ɓ�ҜbyJs��?��v�"K����2����fʾȦ�8�X��b䣼4���#�"�(Q�"S�r���X�`ɫ�7�,�w�u�h��� 8|���H���F�)%WH�!���� RU�P	{  TIn�¹�N# 	QɅrE*�kVQ3M̤s�A�j��HsD��IC4�6xb�3�A}T�`�fO"�N����F�n�U�p��斃��H&h0��;
��<G$���5;�23�č�7
�ɼ��kU��y��F������*3،YrΩ0��0��E@+&�Vۆ��ɂ	�ĴTZ��32wv�ѲW�]t'&עx��̉�b`w��C`�p&���d)	4�D�j�n8�9l�T&[e7���D��=��%'XN� ��hRf�^eY%Ǟ��{wGUU+�Q?�ے�/�wDhL ��u-��	 �p����#�yIrt*!q7XߦJx�"���T�( Y�����/$�
�1���?�c�"�9
YY�VK8�xpi�ɶT�B���)d�Q�-U�Ổ3��~�����BX���!猜�{Z�VT9���ѳ�~��po�^U��OwG��^�#�  �䅺y�_T��(��̑�r6�	B�Q!%�dk��f����u��W��s�YS��Y�3��[/6��Q��"}W���G#y�g?3ܼ�_��߿0r�w&�%�z�/���^����o{G��cכS�>�jJ�> LsG6I�yD�q"��J�} [  _tc�0w9�\']��9B�DHt�ف{�.k8O
�#�$�$�����] �ٲ���M�?� Ě�ݕ܌:�	�z�P�t�v1�aQL{F�ܤ��~���9S�W0�\U�8qq���. ��� n��+7ew'rnĮV;�ʈ�027�I�9� ��X��lv��~���f^���5��D���>H�>r/�WNNH�N`�5n֐#j�v���LD�w*�+rSm�Zkֱ�n��&���	d�bV-�h��Z/3���݋�X�HD�� D]���̹�W�݃����:w��9�����Lp��^�A�A���;�ɉظ /Vբi�kp�`���(ʒ�����'DH)���w�O��-KϚY�T{�a��B�{Ť`��7L�,+�:V@1��RiԠ�W��������3��$>"Z'�Ĳ�I\�X,���DTHM��b�0� �ݠ�@�7K�k DG߇nI�j�@D� �z̡��H!J�<'�d�)�Ua�����~�	q_�=�	N�����B���Z���C�ê9���K̣+fU@���'kǮG�1�x���`.���'���\�4f�۶(��yE��e�����N{I�<�������c���!Z�3\��3/`�U����b�:�(�Q���X�3���;��z&vx8�=�y�鄾w���<�l�A�O�#\�*����y ���$�b
 l1r�NA��F��Rm�L3yUQ��r�1��R��*5J�Q��:��SͰ�������H0{K\���8�{�F�L[IiˍX	yf��2���p##�A<� V��=O�hDN� �-�_��TGL��Da���;^�=3sΑ,o�c�=m�9���0� �+Sq'*N?%�s"	3�q6��W�:�[e�FnV�Y�Z݈X�qK���qf�� �������� g�VnV�i�����;@�O��DJLF��ff�e���4�p h����Ǡ�Tw6w�AV w_y�/e�����߯�R(�G���į�8jc��o�-��1FQ/jUOO�W�K:�
+��)P��#�  ���K��o�R�)�$a���$���8���ă԰�yL|��	���j�Q���ĝ~��k>�7VIV*��Cv:ξ�b�\=��,GJN_�J���Y�����R~��{�p?�z���'{�Ҥ=��} ��'="q'�8p��=���B9(���A�z;)=P�$����7O�8�p��u�]�����<����POƷ�i�|��v)��໢~7v#����?>W6�L�&}/~�7'�}�ߚ_��[�ίx��&u�'��nF#v4��0	��]�Φ���6f0�=��� 8��8$Np"U�"�)�m1s���%&f%|�@���u��P�fp�LN�`��Y��j}�J Nŗ�j��Ld)�F�1���C ����t0�N���U@�wJ�ٜ�H�wg7��������{/�2���SQ���c�Y�Y��ưB��Fn&�ΰ��Dȣ��+R?S���/�Xg��8��RQ�nK����v�� C�W�C�ɒ�D�_�ލ݀�����,e��� �z̄�z��������V
�Mv�o0	�lP3�X��٬�f>V���=���|�oR�9H�?^��ޠ�4v�p�$�H�2i�������K��c�ԣ���,�dk��_O�ζ���okHǺ�����{$0N'C[���ܩ�ޞ����>K���pd�]U������I?Y*���[8����pc8�5�F`éF�lc�X@I�!̺�EB���p�;c�� �8���[����o��)N�^�����jvv��o'��v8��g��1"�L���Cĩ۟o33�#S!x2*
���($�̂�I�/����
+��Ɉ( 'b#"��<�*͹���dfK���`��o�ۑBS���(RE��?���BÛ��3p.��y;��2�����j11X�L_�ļ<^�BsK	q���������K?U]�9�<�99�嚭?����Z��В��1I�8YS\����f2�Q1��Tw��k>S�2�/���p������P[�A#�\W��-o31�m_�>N�xP��I��0H��'f����VHn)Kލ�H�~ߓ״����u��	F<��~l��G��u���={�ZR��|vm@��i?�|���jWʓ�����Ǖ�ӈߙ��`���-�bZ?��wZ�����~;��BO�N)A	�!}�ZL����@4�*R�Xd�֣�k&�;K[/c{��!ϧʹ��ǿ����`m�m��a��ʕ+�W^�V���7*������~��`ވD mآ��lPYV��l��T[��ӑ��ia+�F�<$ ĸ$; V�8��t��V�&mf0�š��b��Ӿ'Ho#�S���IA. {o�Q��۝A'�*F��t">Rݖ�G�h���ݱS5`+oĞ�e �� ��0�2�9JTa��&ͶT�Ыi0�3 ��5��2�r/��i���i���v���
�^�0�ș��i
��Q�{�nu���W�_U��O�A�r�A������]�OW0_�n=Ni+�`�S2F�����x<�w������jI>9��k��s�YVR�<�yW=߷ߐb夯�i��)\�|Y���*J�����5J�Z���g]I�v�ώ�[�BBP�U��z�������Pwp3�����nF��ۉ�;�lr'�r��o����T6���T�^���t��֔��M�e����<G$�N��en��];C�4ݛ����+����+���g���:�)��8d�8�J	�2����8�s�����L, J�'�P��86�y?Xi�X��i�{�� �B��p�\��J�C��T�ݏ�5+��I_0 �37���6�,� (�w�lH�� �^a��|٧�  ʺt�&/�E�bf,zG����������~�tr���}߭:���!���'�=Y�>��`�Y-��C}*<���SQǎ���)���>?p����q-�u���>P�}�`�U��)��ʳ=��W�>j���B��o�����K�?�D����K^s~[�~ZS=��~@Ik�����71� ���e"��>�al���5Gj����9��(&{��F}��z�0Q4a�?G�b���b,:C��j���4�݄�37:fN�9�����t�
�9����߬_~�VuYh�}=x���E��!��!'CUai"*?|�#�����:KW|� (iQ,��x9^*C�������'/D0:!�����	� �!��2R��p_M����&gD�BV�$w)`}`�����܏���g�c��<~�t_�-���A�S��>q�w@� !�rF)iO�2  �s�{��4���<곤�Ẳ~���~G�vX�!��r2R@��>`���_�{N���QV�J"Z:嗈����X�����'�>��+���K�Ø���K�����$��9
�!��U\����W�e����8�(]k���9?�R���!�]��T�p�Rut���]�m^4�3��5�זkH咉= ���e�=Z�b���!N+�V��P꾟���r����~8�qQ���\y�`���
bU^|�6P�Te2�q����<n��ξ%�e��կ~o�{��]|��L<�x�̻����zwwk2鴍i˃��5����v0kǮ���y��C�Y�E(�Tn���1�ʭ�C�QCZ�..��X9oO�ZH�z.����|eK�B%����0Z��R�A�q����=v����Y�|r{�vi�<P@~���~?�C:�#��Z���)���{U];F�؏)pG�6x�o5�jJ �|�OӀ��o�߸f\!���������    IDAT�$��8�ϱ��ȼt���z����OS?W�'�z�����'�,��`�����a�~������B�\���lҴ��2K��Wa�H�٥�{<�E�.	��~���#z�=�����pߠ�Rڠ�?h;1���e�%Vp��� F@]�`N0� �1�@�����i��P�I�OM�Z������}n����ި~��3D���_���Nr;��h��^|���^�����k�qp��)c2ق�G���Ї�a�~q��Ѥ�:��䬧�� "䜗~|Gj-#�Vsku���;$��$�p�ĺ:���l5��0۲ݫy����$m'ɓ∤�cqL?-I��>,1���պ��|�uߵ���6�"�Q*N>�m���A�?|�S����m�R�c�5s���g��a��q닝��܁O���엎���|��%�{��u)O�<�8 ��9�C���}���x����֚�g?߶������� 60)�2� ����Pw�W�8��$0`��jBA�'u�C!����p0N���}p��� �!���o��k�(.���H�9����`q�+�Ҵm�'?EY�F"��{�=�p�nE�s��9c�"N
�`\J��}���&���������3��úIeݠ�I�yI�:���y���4Y�'�,>_]��u���دo���?����>z��mI�J�w�X�Dq{ƶ�?���K�i��*!Lq��tuK�?�P����0S��������n��o���ݟ�4��;� G�*���V_W_ކr1�0�DwS=��t��s����"��"h��߿{�֭�ǗO��3Y���ŗ�~���/�Qg��������TY��;Mڶ��8��3�w)Y�w?=���P	'�/M@�O��q��� �Xg"|�����>}R����<�5}��w���d?|�׷w�NN?~�Ԙ�(Ռ>�h��j�<<�'"!,-UU��k4M���QU1�Ǆ&61��
"		���7PI��N}��@(�KAd�H s!��~-�չ�� ������j���֎����*�q�ɖ������9���Έ���_Lo���F�����ة�EWј+{9R�1����·�;<��B�G� "ǖ@Zg�|�<c�ͭ��཯��D�2��F��A�^�}>��Ügu0y�y�{<;��Gy������q���8����X�2Ƈ���@eUA����������R��ޑoq��_�w<۝��
�s+I�ѡ��g���fF�]V���SXv$�% �J �$j��Q�FK׉�����Wz���3>�ן��HmB���l��E
���D��.��ю���9�7[\��\�ݴI���F�._���4[)3�_a���<����T�"�Ï[��V[��*���`K����zp�J�;�ez�#��u)�����I�����bR��O���?��u�����V����������ó�<:
�)k�:�O�>X|Č�nB@UU��
�
&,�8	;��KB}%"\�
�sԁʋ�;̙ �LMܝ��9�,-/s�dG�Nd�rMc��7��c���sAoI꯯���}��yI|sF���6��yֹucS��"�#�c�x�vƷ�`��	��,�'}׮	�_���[ �mH�F��ۃ�����ѭ�؇uC��R�;���;(��2������qz�+eyC%�r�9K�{R��*�|p2��4���a�ϯ��X!|�#ĒŬ�i!5��k���T�-H�8�D�2�1�q�T���"sr'"cH�E���%_1�G0�Y͂U���!��S]J<d'�`���,�D�S�/h�XFk��y�L���� kA!T�b*]�9������,�����`�{/�7���?X�U|�O5>R��+W��Wn�F����	o��z�s;��������l7�L�@���f�$|�
�O��9ͻ}:�eb���b��WV�~�C��*���M�q��I������I7�=m|܁�h�Q߯���x@�>�����r�֑�cfNT�B���	������������q����B�ma!̉E2�nj�Djf�UM-#e����]ۉjY�@�ܞL�D�����*檪�X���bfFo����^�t`u�l)���ݾ�Mj|>�g�,��U%x��@nI+&e��]���i-�+_����5k n�i�GD����_U����2���T[����?�n�w�޾��f��2X#�t�-|x�'a�%�F�jC�MF���� ��{q����sr����r�=��p���"~��?N��iWK���}�����G9�3��w��������n����W����Fy�>���c�d�`:ckk�QS�:ƅHh�� �j�9+���������fN9!���Y6�dj9gqgu3/Q�啟lC�Pa�����2sF���AU�,B�N}ri���,��,=]V"��Ւ?\��m����zOЬU�d�� u�!�6g��Q����^y�[���ؘy?�x���+W����V��ua2B�������t���������9	�W�_>��sFJ	A�N��t,��1��P��J2cC?8�01�oOg�|���'}ܳ�I�78����5|^X>
�>��ݫ}Gc�t�U"oG���4�$	�� �W735SS�;����)�T3g$r,�mx� c"���%rd��ȍ9���� �  �3S`��Zq��@U��s�4U誶3tI�@�'�a(�C�ə�劉}�V��� ��VҘe#�T�����dg���>4���D�ݽ[��gOqd�&_��_��\�_���1�zȵՠ��ٝ������c��R:��w0�����
�y/��.'8;�* \��J0����|�n��r.�idYY�#3��Z�+H�ݔ�PZλ}��yq5��<i'`}����~;���i�_���i���y�i�uJ��Nj�۾u.�O2�H�^R�ر��"��7l�jL&4�������%p���	��[#fN #��	� _U�7�5= ���vx+ �|DBu�p�1��Y����تCU[j_��4� �Ч���*
��qN9�9�)�kS<�/0o3�ڤ��� 3LE�vƎR�6f�ˎP��XCUP��Cr��A�x8j�w.=�'Jp%��o6�_6��N�C`o~������3��������"vQI�y�/՘����蕶;����V{0����)��� ���fĩC�������u�瞿�K�.a:�b6�������w�.�Z����~zr���,89��~^]x���6���bu��~�U���fAU���5B]�V71��SA�ٲiVPb�d$���C�]��D��s�w��]�n�����s�������� �v�����?���k�x�G�ɔȦ��9���5@� "����R6�='!"&�:�ZוrS��Lc'�!d��?9 �e�P��8�7�, ��5L�բ�	b�ȠI�"�L�*3`���܅�����)<i��_�����6�9F��ط���]��^�ŝ�Xg��1?����K��]Y�k�,=���Tu�[Q���f���~�~/�������������],�8Β4:֮U�)y4���rR���n��''�#�{i3- ,�QSa<��:��d���]���)�Y��V�_w)�����_(�w�!����Y��?���iFYj���Kӗ���3��a�ۉ~�7S�������}��H��=m�N��*[�:����/��9���McbrS07ĸ��dA���-;)H��'�]�$V�;�Go�-���(��()窊�0������bz݉G��ҿ:����'I��K_�&u�c;a1�)�4�2��^�D/���7ݻ��.u]/#tO��V�݃�y��䏙��(I�U=ťK���W�u���..=?��d
!�Çڡ]d�ԏ��A�;��s� ��i��6�pޜ�R9!@�4>]�=�ow��g>z�x֯o���#j�'O��a�op��� *)�����4�WU�	�"��H��J�� 㞃�5���?���)�Jh��q���X/|��<�ߞ�m��u���g:�N�ƍ�����ڵk����T���!u8�����O��>�į0���>�S�m�6����B�,�w&�ö����:�_hZ	�x�~_�	�}(L�M�$��PW�Uu%�źr�W]����ՐfѶ�	��≑�˗/ǪJ�h�O����\�ؾ���Wg�����/�j#��k�e Ūo��7�i�w	N@
�x�X&P�����jR��C�w�{��-��a� [��4����ն~�m>9	��g�7,�4�PUT̌�|��_�w�>�89�G�_y�+/s��59��s"����:'�@|/�����2�7�����\U�J����W! \U6��Ӆ� pJ[���<���oܸ�� �7�x�oݺE�/_�7�dŽ�_�v́��ۋ�sU�D���������_��k��M^��?�.χ�_c�_�L}������Ȗ���XJ2?,��@��F�����S�V�gAq�����8U�(ֱ�+a���+�w�t�]0���+���� �T�z�ˣ�횦��4����(��������ˇ��/T�
A"rJМ� �Ӄ4��qe�|�f�%|�N�!�1�z���Ӌ�nM����* �	)`1���|��v=�u ��x$��9�V��y�� ���OK�1(|��[[[����|9�e�σ��qj|܁Ow �:�W�{ځROkۿ���x�OWD"��H0OP�U�U�@�ݡ����3�����ڬ`����������ٍ~��^��R]�	���,�(�5��trX����4�F|�+_�����o����bs����{W._�������ƍ �/_0q]���_��=UM/���sq�"�����O�v5���:�QMG]ʵ�s���3sf"g@f
�$>��a �%�,$%P��!"�5ƓI[ג��S�uf�����J4����������-�%<�w�ʕ�4V��Ӧ��RK���-�����K9�q]���03��s03�FJ���3�z�7�)A���8ߠ˜a� � j"�"�d%<w�yT�B�D����A8!�C���T;ޣ���?���u���?����^�F�P���mۢm��ҏ*��Ӟ�?��i�_���9�����������=����5r���*�'%8+1w!63�|Й�:�/�eN򝪵?�������/��k4�ϫ�~������b�@�Q�9���Q��㺙T�d�ĉ��gf���Z4�{��s�����ޞ���/_��/��������������/��a�ʡ5�f�R7�@{ �CgPG����+�Bdf��vPSD$
��㣌�Ď�$]@VI ��q��*����HB ��kSp�Y��W^��t6��͛77��3�'B�&�I|^���V]�"��|v��pߩ뚘�Ѷ-��1��l6�0�L��\q��Wp^ҧp' �5�"����h�!����q�x$ :�3��[3��6<K���i���>�n5��d4���z����������=���=�'�t<����񒾓/t@I�B@�IH�,1	s���~� ���?0�n��>�����ʅш�����l63`��u-�k"��@3��0�ɸ�Z�!��
&NW"�$�:�h�9�d2�w�y��|�M�|�2-�L&��/����� �����o;���޾���Q]��� �Ax?V��l�97�5V�� b ��\-2-鼺sN�D� p��8�����V7�k���J�����[��ao{���×�Z,���9>cx��~��~����1}>��_U�WB75-�/�/��@�BN����7y�,9�;�fo�%��̬\j�D���dG��Ü�0#s ��SꯘO�r���#S�&��!d�[�=+��×�����y�gT�R�,�����#��m��}���jl�ꉦ�K���&�1W�8�ZTŐ�\~Y��Q)PM�u S]{����,"n����2&V#��6�r�%��.��]&�]��QTJ�Ή)PWC����nd$��"��su�6xR��c]���\93#Ɯ��,K�?[�EO�Yz�΅�w1I,Hߢ�岥�v;�:~�+�q�h����<Q~M���Y*ۋ^��B=��̞�}�=���X�w%
�v�����%�v�ųr�˞�����Ҿ����{��O>��%;��by {�����%���E�i�?��?��@K�����-O�QR���H��tx/�W+�+U¨+�ՙ��KE
���_�ݏ�[���t<�:쿴9���ɿ���_������+>��Ѝ|c�@k���S�2UfV�5X4$E!�h`S@C���A�3���,�=��g�{�=��?�g<x�@���x��!�o��?�) K �ө��_���W�������<)�� �w�ӥBLDER�O*t��#!�H�ǻ@̵{�#	o���pf�D�%,u�)\IJ
�����(���r6D��HrZݼ��&�ϤM?�X?��%����X����˕�~8�x���E廱�7ۮ'�.��B& �W���D��D����50-)�cN%S
��_@����ӆ�٬!�D2!%#�\�1Gg	}1ƥ������:�����UbA��[��[rGRۉ�}M��u���ܟ�F�ğu�g���'������/�ٺ�P?�{�>DdA#�iۯ/�^�1��<}�_�<��~��Χ)�2��倫�TQ���pYԃ*y�A(�>�r�D�؝t������D}X9;�"���r��Ϳiy/w��`௪��"U��R����
s��`f1�yT���ټ��ҹ��UA]��VA��Q5gÿ���2���{v��m>���Nj�ш۷o��۷�ʕ+:��h4���?o��"�,����R�w���'j&�L��BũvmG�h/���q��0lH_��l���)$�/�IA�W�F�4ճA]I=(�:_t��d�KH���\�t4��}��¢w0�Bw�B��l`!�E��2x�y���G~�H�耖���!-R��z�2R3���|�5�7�"ZҴ�vi��ug$b<w��J}s�Χ�Yv� �d�_��"Wy��4MKJ��)�|��_�Ó��Y��I�+/���� �.|��=ksu]RxD�s޷��M����[���ck?�+{����z$�f�SR������ӔJBU�eт�"&�m��Sl�R�M:��������������ߗ�÷������EU)�g�B�`�y�y�=tg�}=9�& ��]�����דɤ�'':�yY��ʪtq�EIm���w�N܉+$,qJ�̈́�KOȨbNI_|�RL��������*� �lg�}���}�/�B���:��0��"�(�T`H��,&qy���f�	y��b���8j�D��'�����{w?e0t�*��`c{D]�ܸ�&�yG�%��I��LL�I$�qX&{�Ƚ�ҩ����fvj�[�vAϓ�K\��F�k�?�\�������W������8_cvA�ʲ�����w"�9W�!Y0ѓ$|<����%~��do8�ι�?��4��I�O.�$e�K�Ue�4�YJqn1��Kݏ�ſ,����4����O�@x�w�w���n������M&p��������4�`�B��/��q��b[&�J��ŅXk3���tFJm��U�ˀ�����L=�o���}�YP�d���P%�����v�Νˇ��B���@uh�%+���>S��0�I�R�\����_�{WLs�Lb���`�i���wLg�|����XU��
W����u�̛�d�2o~�����
e1rZxmlp: �w��y�ނ�-��2��]`Q��-�2������l8��л�W�����$K��ئ��EMQID;�4$$$�6L�毛��/���;W�p6Ҵ2��h�r�i ݊�t��u�d��*T]���.���nA������� ����ߓ��=K>��]93��F�k�ʂ(�֩�#1)}�����fBe!�Z����D/�-�������ԏ���	d��B��묒��=    IDATj
�����%~o�"H�Tf� �@x���8������'��'w�G\~}/�mrܽh�E eل����!%v�fT�x���Y_��S�V
VV7�q3qp8�`�������]��Uw�#��	~� ,�<_t/[/.�Ó��M�|ON�l���}A���,}����x�{����eq߽�e��"��!."�d�����>�7�_:;�����:�IUuiY�~�e���(��Ƶ����n��E�я`��+{�'L���hu�b���9��]<��M�Mև�+���z=F��;�R]U�h4�)��e�Y��S�ŔT�,�ixt�\�Ϟ[13�>h�""`q^J<��[���x1�]�:D�h�>�-O��,}O�$�����D�.�jUI6�R
�����1�W���HUU�llq�֫<x𐽃�>RՈ]`y@�&R��ћ���� �ǉ������$8�:�����*�|����-}$�����,Q�9)�Fq>����ʹ���tP��u-�9��,'[U��%1��AV'���7:޹����v�������;X-�0����ae��}_���Ͻğ�����m�d+��j6�B5/g�]ȁݽw�=v�x��]H����0��RBP3K*�daݻ|��x��'`s睈8�d�X�3�>�����$!�"��\GY@�L�{��~�)��̍y����u��+����d82�#�M{�."|˯ǥ'9M)���ey�����%~��h.�b�u=�^3�)����R��y�m��]���ڞ����i~ûr�T���Ih���������	�N]�-��Ģ(���l��?���pؑ>��7�~��"�9�J�5x'V�SAI�"��;���v^���B���B����bT�G_I�\��/$e˛7w*_��\�uD^�m�>�M�'�$�47���I��`�9Y�x�;pa2?M9!��֧QE���"�*9�`��%���
�j�`8,&�M3crrL�-�tc])\AQ��m����nҋ�$����h/��-o�eqQ�/���c.�^��E�]��,iXvO^�%|Z_[>��sXN*������'eٲs�<����{s���y�e�ڦ_7����Г��Y������N�~�۩#�<���+��K�Խ����}R�vP��	�!bw$���l��]4x'�t큨�aR
W���b{o8l���w�?�����-�?��]�r%m\ۈι���w��^��~P��4�:�𾬮�q�bW�a*"&��oڎ�sڕ�
�����{"���
�AL�}E4�dB4c4�`XNU˪t&�"El�0��7ҹ�����r���ⅸw���
��c�0Srֻ���/�v[�&:���>tP(ԑĐZT<b��N9<إ���R�c��7�׹r�%f�#�r|�K��B>�CBw:q���m�8Q�yvY�.��N�[J�4�vY+vѤ��-_���C_��t_�-�c�"�:X�D�@41|մ)>��O��^Ǽ��8�bU%G�,��jw����oۯ����^ 1ѽ������y`S������λ�
����QxM�sVz��� G�Fy4��4M����)K�)�H��,��Kf��@;�L��%�h�b4}�w�ŋ��L�,��">�[�I�����J�)���)��=�D��S���L��y�����G�mlqu{���m,�f���N�ɹ���.�}�O"/�-���r$��g��2ֈ��w>P���w�|�c>+.J��~Z����/p�2��%ΐD��X���d�]A�Pj�k�4�s1��hP=����]�[Yv�FGP�JU%��`.��Kkc��������o	_ j� X
�6��G�?U�êPV�P͊b:oO=O�պC��9�>y{��yz���!D��d2�L����j�r�r��"X���P��h��1�S�p��]|��|�JD=Ε�#E!�4�f����'���������{|���?�'����ō7�y�:u]�
f����O%ςǹD/
t�Ȣ�8·��������$�����R�|U��ǹ���:^���%�E����Z�5N���T}0\4��G�(E��$wp�uM�s�jʔbi�v�4���_����H��B���h2(��{T��)�#�bJI��[Y��**�f�)W�z���AEL%��=+]�	X�	�������5���g����=qV��ʤ����d�u����a�ڳ��jf�tB��Z��C<%��, )�.��HsT$'�4GJs�'�����U�Xl�������k|��B;�0�6�F����N�9*��`�(=Ɠ4\O��=O��]Tw!����=.j�q�b��|��'E_��T�=g�����]�d�T����Lܤ�⯕�~�CZk��%on�������{��?��Ye�nؾ��_���o[�/�/�#W��;'���ʪ�(�<�R/7gɥ����ޣ3d��q*�T0�f����r���ݻ���e5,j�J�����f_b��~l��p���*�{BLfǄ��5�;�־�˱�F�"1u��M�
�D�3��y�{���}�\Y�� "�F#����z�*��Cf����J�mp�u�l�Zvc�6ھq~�͜��ҷ����/�z�h:���z�o/r__��t\�M^,����p.�iJ�rb�U-�|!)kG1�4�Y%���龰�?p���h���߯Zw�?����R]��
@<f�qP�n�L�!K����c&���z��㜊�Unv�N��a�I�k��0<7�[��TW�1&�����$���x<��_�֭[E�d2�������5=Yr9�X$u��라9� �, �9>�����GL&ڕ��,����ƍ<������,J~1��H�����:���"��eH�E�E�_&Z�����/Z۷x_�h|�=X��oï��^�(��C�ab9%HNπz�	�D��Ĕ,&u]w��/Z5_�pD�/
k6�7����i|ݸ>
+��mU���B����[)���,��e��v��4������=Yg��91��/�y��L���HU�n��;�\�o ���5]�E��5��1���ƾV�eI�u������ܾ}���888���K���%���:	�D�����J�ZrTՀ��rxx�����'��+���:����F#�s�S��d��e�ȹek߂�<k���n�/�'���i��ߕ��|���1O�fa�\��"��R�w�K,����ɢE_�����M'|>p铨j�-K�$�Ɖ�WW>�����VnnŮ���V��;gj&�E�s�[�
�h�o;�,*�8�w✊����RS*����ߗw�yǿ��;�Qx�?</��
ZO�f�%M�S�^L��Y���U!����^	�0H��#+M�� �Rp�"�W���8�5�l��}dJ�njC���ʛ���K�)7ߒ	Ww����������x�QY�U�æ#T�(Ig�2�Ѯ�3\���-���:��G||?�ze���IG7����u�+N�#�UX��CB�����(��$�|͋6YT�(��&8�)6��QB��9ae4 !�.��Ɣ�*�2��]G�W�$�	)���dXה*��Z�%|YR�
N)�m�41�LH� BhI��f��Afm0��7D�1��x�D�xQ]�]�=B��GB	(�(f���U5�@�em�fm͑bK�[�V`]��(E�h��pP���`�����ONh�Hj]H!2�$���%�0�Zʲ����|�&|m����nѻ{W|o�}=M;��ܻ�y�ߚ����Q�v���� G�bN����<��L�E�'��FD"��E^T��� uG��w�ύh��&��P�[�-d+jjs�V�9��l��ǜ�R����I�eH��hF�Pf��b�!֟B��GBBp�ߵ�v}PB����Ғ!��G�C��1E�A]��<��N��
�\�H\��b�1:�m�B𑤑 "������.�,�GI��Hj$I�CA۶e	>��Dт.��%j�R��@U1͙�N��k�x�b��༼a���J©�Ԑ�0u6�4���F�릙+�L�a��o����{��J��6�\�t?|�*J�K����_����˓�ͦ��n��5�BKW���T�y2T���H1��D�{�-Ɖlau���9�'�6��>tz�ʊI�Z�|��W�ջԑ�������Gw���:��_^Hʖ�$�r�y���V�%��$�rF۹��Ia���R캆v�B`8T�j��W^e}m1��>��#&�-P4E����B�����4���ܿw��W�P;�Kc0������&m�f�'yB{��X��-/�c��J�B�������Q�pP�:�4����l�t2�x:cg�hF	\]Ǥ4M��guu���5��֩
�w��}�����g�]���.$�]������L�)"1�$e�Or�*/ζwV���b��9�$W����v���u}����eX�z��8:�Ӷ0���!����9�`�>�~�!~�v�?@D�q����ҮO ngD]EP[��G���;l���rf�,�>#������qQ�_tϟ���CDR�$���b��0�$ 2q��dFgж-��E�c� ER��cR���dK��"��9M�[pYV�1&F�F�Gj(j$�#.�G �tr�^�!��������m���yҢ���_�����'�X(Y�H��9�-�B�RD5"^Q�UE�HRC\n�$	R��8<"�� �)R���S
W���fGQ�"���=J)1�:,����:O��̗5���Ec��gfQ̢z�$1o�pH�vʣ*s�L�=t?����}a'���!��M�lX�8�9y�R��=[s�%<�<�,�$b����s"�D�j�hf)��߿.�o��{��?������GL��������eaQF���=v�>U�r)3�'�$�+�	0��d2���{�ܿ��X_�Yٹ�p���gv�p|<e2��"u]0K1[eW�z�	�D� "�63�����2�W���*+�5�_����[L�S���l9Gz���T,��\UYor��67�X�\�\gme��.k 1��89:���]>��3�|�9�Ʉ�:,��Jԕ���1�p��k���k�z�ò�,�{ۗ�h��+�)���@�6��������������w�����w��	�,���O�(��V�^L��Kp����-����[ߺ�͗6Y]U,uЖ�d:�<��Ǭ���o����xX�K'�����9���h�"ބz�M����H�^�Ef�D���8=	����蟉�2AL=�9�0�����:�D�[E���\Љ��D/ƗɞWn	���l���?��	ƫ�|��
������&���J�D��t��p�Zb�������r*�̄����5������e�C�D4!�e�-9�f�)[��`���Y-%0��zo�|!����f*�rZ&�����4�u��Ήa* ��G��>�g/�W���p���DOz�]�L1��s��O���m�SB8ˉ��@"�U]`�ֻe߳����8�""�Du&��P��+dg>E�೎/���ƻ��������_�8�MD$���3U��~���X�N�I$��&̒8����Ԉ9�yդ�h2�����:�o�?z��O�n��Ē�9AΖ�_�b՜�(5�I�G���ߣ�;��"tDli��(|�O&G|��8_҄�nMp~���5��<b��>'�S&��m�fWMO��'}Q<N��f)[v��޿�gkk\���K;#�;W_��˯p��}��'��UD����b�]��k�����׾�[o���[��X��RQy�I�*
�ʓB�l�p���hQrr<a:��R���Q��Q�%W��������;�e{c�A�
ɒm���J�D��хDg�:������m�{�3>�U��;w�����s�e��E�w�U*��>U��A��p�[7_�;����z�����)6İJU�����.
?�iM���g<Nܺ�&��X[����s>��
'�m�	�*N ��}A�	�ق�-89�֩����I�)���]�w6񞒼Ǻ̗�\�*zRG�\m�@�X�/�u�ؿgbɤNL!H��M:{�Eu�t}�29���"!�P'x)p^Q�ݜ�v����]����M|?��߱�6_�إ����1g�i�3�xvOK�{9�5d]G" >���؞�W�!����Tɦ�6Sn�9��Ϸ�'��9���{�$/`�?�GWdKe"��ĮG#�@��|%�-��BL	'�� a��.y�5�O�ED��&��,!Qi���Hw�n��YbE��1�����:�Ǣ�vU�C�}pN������2@_����Bԩ�:ˉ���W�G���.�|�0�K�EM��>g3�#Q����$�ߥŔ�����8=���σ!�pb4�)w�|B�ɢ(����aUS�6ؾ�
/�v�|�§qxrHA�a[�i4��EOnP�	��|:a����L�W�յ-��t���)�=d�Ͳ�/٩��qH)���S��<U�,K���x�����w�ŭ��3('���$u���']���������](IB�y��5������׹v�5���Qj�e�DBgFH�������kEQ��oP���ؠ��/����R�k�Ǔ-��5����^ӂ�H�=�p��K��\���t�	�k�h�������6��P-UA:
/x�Yۺ�`4�HI���=�yC"���;�uH!���N?�O�-2�ҩ<�{.+٪y���Gc���v��[-��M�������!�d�����uvCg��ٓ,��P�:��@�ԏ1[�]�O�ʧ&QA{k�j&��소)[������W�=�_\vz�2Ձw�ښR"Z������T��-�Kz�Z"�EW��j-���RB,��e)e�j2�E�1eˍ�C]�J&X�Zx::��� �9!u${H2�Σa�A+h�Ę�EYP��y�h�/�+=E�yAd)�6�4�K�b��H�w2>��-0���߈�L͂!��ⱘ��W�Y-���o���i��&bD$?7jΝe]83�\���4]�Vg�R����{s��z/�S�n�0uw�|c\��x1e�4&�E fk��<��w�pI��+l!8�~�]ly���3I��C������b2f�������JO��-v6j�шՍk�|�!v��m�MNH*$K��\����(��YJ��b��落�����2�`<������5��'Nf�E�.,��E�Lr{g��pu�j��jM#Ncv�i��󖮝�4{w9>>f��h�&뵊Q��($E9b0�`P���D-�fmG;��t%X�F�o�h��y��0ZYa0,����2�]��|���!���]�/9\|��Mx0���b�e�/kB�bN�ݵ����>L�S��GH���56�����Wj�VG���
�+�ll�ě������O~�t:�=>A,�4�-N-����
��ɹ���'�D>�@��h�x�כ�Xv���]Om5���GJ�.�g��D9d8K�9uX�P�M�Z.����s�E�Qu�k˚y����8�p�'���2��|�!e͞�~��k?S�:����ړ��I2���B,I�X���%�1�]��%��^��\~&GÚ��eRo �Q�\ͧ���-s��U=��=U�y���L�9��	M�е-��u�)����*����>k�����*!VV�X[[��+��$��	M;gz��.[lEN�/�Ӭ}Y�����a�H�%K!�4 �˔$�nv�8�pxX��;u�b�*`�K�_�a�["~}�?5�EQJYV� a�N�N4�>��?|x�)N�K���H��۷=쓒&g��Ÿ���a<�l�[rS�Z��K�I�)�)i3��D�J��a�if�ܻ�	X Ԟ�^��+׮1v��q	��f�C����H@�1��h��I!`��"�9��c������\�2��W�X��a�����C��%�S�ڴ7H��d�G�ޣ��̚�q]��1`\WĶ�d:c���}~�{w�ppp������ߧm��Ρ�A���pEEQV��6U�5S��vyp�{�G4�zw�pr�G�Z�j0b��^�z���V�ͭ���C�2�n&�y�|��FL�l_��hD{7�"�	`JB� ���p��>�����    IDAT�����|�*eI=2����ڕm�]������!��*W���`��������1��N^Յ�,��Y6'8�42TD���)U�yr������%F��E�ʙ'HUz헜Z�R���αUQa���"��k�򂤯� �KS��Q�1s��(}EU8W�
Ż�d�')v�d���ު���j�Eژ�UU�����0��c ����5�vJhbꭔ�E�`KOZ�wc��Ĥ9��N��/D���^�[��VB����sTUE]E��8<4��	)�)�(r_Ԓ.u�%k�o�2���w����l����|�	��1 �0R�'�]��<�������+�5��ܽ��'�E�h8fc�7n������늢�E&�C����}��qpp�H"���/�%W�!j�,�!�R�
# �Q�>~&^�Ǉ� IUI4�L>�"`@]�Rץ��Z#!&	M(�s�{��B1��i[�Yx.�W׵��t�%"9�o������:��{g��lh_�J�'61��B�@�k"Ė���Ķ�XK,
��`m��z����:x���]<���fKR#Y�cy�.��L:,�ل��#hژ����5�zؓ�D�F��vq��u�#n^��:NNN���A�uL�'ܸ����q�����������_���l�rT�s�e���W�!�+�,�e�#�4͌�Ç|����/~�ǟ��d��FO2!t]H���V7���-fM�q�Ǭ�\y���s��O��ϘL���~���ˡ'B�~�(&S�	E&$�&����?�o�����ܶs���yO{��+�U�W�\�Wn����o����:�(hlll0��S5���XZL��w��&�����}x�4��ʗ��_�,t�
KZP�>PDZI�������G�ѣi�k�"!5���Ɩ�����ら�~�>��f���ˬ�����J=P�5E]�R�ifL&�̧��9�����v6��|]�Țؔ���pȵk7x������u�
];ez|���}��a��=��t˜�}!	E֪�Հ��-����rt����=fwwYT�[�Bz�bo&	⠨+VWW������:+�1�~����9��4�H����Sams���|���x��ׯ1��������)���D��'|��'�u�g�9xpb�R���Ң�%h�˯���o��������&�̻@UUl�o�g�����op���S���ݽǝ�?�����l����%s9���pj� Щ���If��c��I���������P\��E�W"-{���A~9�i`�eY�`P�JS�� A�%)���mu���7���e��o������ruSuE,�I2Ra�Y�{1�	�����V��}.D� �]?�)�T��Cb_%aq�G��	]B�H$�w$1b�'���=>��R�z�7^c}|���d��u^y�u������4�)�ù�^����;ʅ�.JW`��	��s%��p��ع������.,�G���<t���eA��u]����;�;����w�bu�fex��h:���G1�Lr����X�R4[L4".��������T>���~�7��_��g��bT4���E�1A�2k#�.��p���m��/��@�������6e�畓�%C�z��/�<a���E BE�T���b8K�4�l�U�"t�޷��<� �I@H���!U5�ƭ[4m��kTU}Z?x:� �SV�m�z�TՀ��b42��ٺ��;9��,�I1�5-��CN���6R����1u=d8Z���fY]]�I�C�����u���(KO]ק�O�L�\��V�ϧt�c�������9:�2�wT��s�S/��W7����3^Y����6k�EAQUT��tQb����{����������î��ҧ{	8�qEE�����o�������IUK��h���}����w�����#U`���D|r���Y�R�cF+�������}���u>��~�ӿ㓓�e���^K�������tμm�Z�d��	�x������笭���l�K&�����pER-!� _���ş���?���q��k+���ks��<m2�YIkc��dkm�O~3��_���kW��!�9�lmo�}�*߽�=��G��@�[7o��+o�֛�amm����ϧ$K�c���Nloƽ{�N����B��������kO4V��;��73�RR����peݚ;��O�#N��$���"2J$ĬO1d��sc�Rt�-��>P�(�Sw$VV%1F��EYX5���j!]�X��R�?wItu�&���[�_'���omŭ�s1r,$�&/�b�­)�q�.+�-m�xߧ49WbLU)ʬ�S���LC�!D�)�n���]�ݽ�����J�)c�\��ε�q���w������k��EB��}^��m98�P��A�+��U9���������a��:����	����f�>�ri� X�t��]/\��f'�A��d�1ϑ�d+'��&�Z2��f8'�pr2���8Ga�� ��8�ݯf����b�{�hh(���Y��3(+�Fe�ꜘ:��J������c2mh�H4��թ�T]q�7��M@�*����֭[\�v���uU}J@;�m|�O��g�?|�g���?c�y��!Z��$aD�V��4������6���:o��W�]cu<ƕIF��S�8��8�EQK̛Yւ����|���_�ɤ��<�/36Gk���k���M�������M����w�:e��x}���Y������ۇ�g�~�����LF�x���Y]]gck���+�olc�cPy��ʠbmu���;|���3�?�Pl�p�hA=�}�*W�^ge}L�"&�ٝ;4M�l�҂�(]�D��`D#�a.��������7YPU>����8�/*:�62�޹���w����׮]a4�4G)�FN=Ml��A<�H�x_CK��-��1{{{Lf-]�9Q��(����D5!�`gg��������_ccm��x��`p��s��Bb6k������=<x�l6���RP��=B���9<�=�>I�)Q3Įn�)�������D����%�8,X���{���B�^��x�$X����������Xx.����8��z3�s�d�l�=z�B�Xʶ�b�E�OK��s[�؄>|��L�'���w5����m6��E�0���]�T5�w�re{�c��Wo��ko�M��p���r`h�R�H�esz��R�tm�d2co����u����YY�dee��f�<�i�����?K�v�09f�	]�S�(r�F\��,��J��>��"@f�,fk\�!��9E��IR������0U���9�MV���˝	����>)j�OA���m$�
�E'BUЀ����� ���,P�!A9j���n��bEYgW�z\�H��h��ԣ1/]���[����os����1������)*_P�R��5�?����
��_����M�����,K�	]H�6ulllp�O�!���?���k�WWr MO2���hq'�z�Eb&{Zd�_j�>8��;�?�Q�
Qq����������z��ׯ�V��AY�Y��5�����@�P�UΏ�uY�N�'��1kZR��S�E���\I��J|5ė�a-lloQ���J�H��u�����mmg��pŀ���y��^��͟���>����R"'=�jf�[;W��wn��[o������~N�3�mnRWbA�r�:߾������W+����4��n��`�(|��y0�:���à�p���������w$s�j�p��xe_V����ޛ,Ir�{~�����1�\��YP @�H^ކ�Lm��`2�B�2Ӫ��3�7��� Z���nKj�� 1՜U��c����8�Y ,Ҭ/�VȪ�ʨH�����N@������p5�V�f:�q9>g>�3[L������S���9:<d>��&	�+N(�p�����^|���/�&(��@Q�����F�sA��������fK�UD��?�m�d�t%:{���xM�<M��tF��s���?O"�v>x�%D|�����*>L��cR�VN��hV1cK�)�=�,��V+�F%,���"6��!K���S�>{-M�;l�;����orvz���*;�#|3~v,��%(DB������t�x��zA�������3jy�?^m��Bo�$��Z΢%�j��뢁��W�|�3K��	��4��� TD���_�Q:�(
�}E���01�!"E�1�g9��+���sͺ��cV����ݨ�B��`��G�C�h�Ӡ�@3&N�,�hM%e]T�QXg��C������;��g��{����W�$x�AI�.��J�f]R�t�nT��NN��0��	(6Z�8�ع�������Oʭ[�h��qL��ZTW�e�"��*�����y�m���ҜCh�r666����w�{�t;�L'E9ie�d�@����0��&K���cgw������\�ˁjQp|z���S���n>���bI��	���k�7TQb�H]+F�9/�/xyrI�u�i������f|9����$1	N��l�D�w��sc��wﰾ��N.��x��K�|���d�B������~�.?�����Z#�R��1GϞr���ň�d�
�BJ�N��dlo�����v6�v��Zo"����fT�RV�����m����~v��z�Y��G����.·L���sF��XE��u��h⬢��O��6]>x-!hq.!H&>t�"7e9��*F?��]�e��e�Y+"b�^y��Kſ���8�Hh솔x	`*�&I^�ܿ��q|�굚�>@AD�	Nh8z�b�����"?��	��&x�m2��5n�챾��.�39=?c>�7#�f�1�V�4����G]MPi�+�<���`���M��6F��m�`��.k�,�b��"7M$��Jc���j泂�tJU
�Q^����������������;�5b�	H�����"c_Or�з�(^V�[E����AB�QT��]���a��G<7(�����a�U;*�s \5�A��A_wQ[5{+�«|��	�ST�F���o+TH1>ڸ�(�A!J�Zy�]���/�.D/�X_�tk�y�������O�m��tp�1��#+���<��ՖD<y�IT���]2��B�E���Ԉ(�����M�~�m~��coo�$m�<,���((˘kt�2:v.`m�s��� �=E9���)O�1�W�J�N����m~����p���<�[Ǽ�y����/�/Jfe�d:��6������:[k=�ַ��V֎���E��
���C|������s��m޸u��A�4Mpa�kT�:��ʯ���WY�$�*���������F> Q���7�����gO(�K��x�#-��������oqcg�V�x...��g_���Cfe�$)e��������wٺ�K�Ip����#>��#?���b�eP��E�v�s{A7ﰵ> ��d-���-�V�Ӌ�_L�$E'm���JR�����ذ-�~������x����,��]��ua��F�%\����~���+|P��H�}Ȕ�\�M�����^zý����s�1~s�ר�\PF<�;'�YQ>i��פ<
(�F7�R���9�	���^_��TP�뵚�?$��/!(V)�MW�'�RE��d���$��u����޽�9ؿ�5�lcΚ,ϥ���J�"�6�F�z�I4�\^����s�n��9�y��.�7vٽ��d6���"*� �K��=7��F�9�x�f��|��)K��G�}fV��W�=V��`S|��-1.N9נs��)�N^N��h��􂁠�C�i�+4����o!�����S�h�5`b�%����EX]^"�P��B�Oy�Z2
\G����H�!&�xoѾ��̅U��M�A��R�G�ΗjL"�VT����=���n߹�;����?a{g�f�(8?�����dBQU�pɀDJ-%��Zl���S:���5(ɘL+T��%�"ow�qc���Gܻw�[wn�j�(���s�<y³g�h�q�S���c�FJ���0"ת�*g\^�svvJQ�h��TB��r��]�}�]���0F���>~ʃGOx��)�Y��(~Q�!�s>�����ҷ�e}='5�4'��D��z���r6gV��rR��]ƣ)�6t;��[x7����ٯp������QB*��$����鈧O�s��.���5�7n�`gs��ጲ��������g��-�N��Y�1Ϗ^���3Ƴ)"-L�Q����6���(C�e�ł�|�pt�x<��/�֓jSq��͠$E�%	"qj��t�����$AJ�$ }v\U�责���9Ϟ<�7��/��8?��\�DE�e���_	/�(�ҳO�`��Q�r�$@)&���BK���y�4|���������g�uxSB���T���[׫�;����%oP%���]Mx��y��������՟��o�X�U&��"�mފ���ky�};�@�]
I${�6��=�֝7IjO+����9NN���8�]fs�k\�
� �����.�y������t�~+es{���999�r4k"IT�͸48$�h�؆=���WYYL&��666�ی�l5Z��(B@y�8�wq̫��#K%t�E$o9b��d(�QhІ�5�ML%E�+t�1LC�F�(�p��Z�H���c��X>D���x���T���W��Wk�<{oc�l��iE�j44���Mu#U1��	E����}��N��`ݜ�Ι/�+��N��������7�bgg�0Ox��9�>���!�јEY`��J6i���@;��{ܻ{���8������9��r�r�hz���͍=~�����~���&y�CUU���~�'���/�#?N����^�ٲn-A�E�ź"�D(Eb4i�����ݻw�qc�ԤX[2�y��1���o9?��|8�v�J[�$A����rD��T6���(���;��+vw�9::��!�@e�x�,j�(n�9�n���D|��Y�_���vH��S��-J�>;"o���;wnq�(v�6������sܼ���0�����}�.7n�@)�t:����|��!�ć�R�� �£Y�Y�{T�o����u�EE(�.M��J���.��798�.����k��D�Ơ���^���΋�>��3~�O����e�yZk�jb݂��]D�}�R�%�k���Z�|[�_w�^{���/���������^6�E�w]e�%H��36ت���X�&K�5��^�h��"���weY�,�V糿�_a�V���tU�:���!z25{�׭���"r��-���`+��Ds~~Ni����Ռ3�`�k�3��(899���)7�{��B��g}s�v;�����j���EH�kޛ֚n�e0�n�ɲ
V�󧨝�|�����B�DH3���z帮>Ռ�B]⛍xxu-��T�Z�(�5X,�ɳ�,K�=�wx�_�����4�n���:_�[>���+�}�k4�$IP!E� ���eFŪ��"tZѤygg���I�YLLg��`��veZnܸ��FDe�G#NNN��ˇ|�駼<:�(
M㥄D�[T��7�����I�#������ޣ�������u�oq�����s���!_|����o9>>FI�l6��Dl���k�)� ����(M��F���^o����v�I���(T���;��Jst�"���9\dI��������&Y#ִJH�k�.F�h���T��J�e�0�/��x��$�#׎�/� �C�L����#=z�����ۨ��	,��^�h��H I2n޼������Q�G�<?<�ɓ'�F#�fZ�(W!:'5i<�"d�6���vsnݺ�Z��%T;��THL�H����kl�]P��H��,Kʲ�A�a�>�G������?棏>�W��Z�h�$*6˸FTuu�,�����]nb���J]�}��u��\KgfM�j������?���~���l�,���[�[7��eL�s�y��^[k��R1Z��t����c�EI\�B��q��R������_|o����z���������tT��G��d    IDAT@�I|���U}�y<�D(M��d�+$�A�����{�TSy�A���Kϋa�f�v�O��ؿ݂`p��#&�)B Q.�?��P�p��ʕx*��0ڒ�0yn8��2�z�<퓦��1;���'�Fl��Ȥ�� m@��.���8&P1] Ҧ.=n1`~vJ���*����7�7�}��W�4�8yV�! ��X�9�c��5�h敥P�"i3��VL�/E�	5$���zM A����$x3��'̫�m��.yk�v��1��$9b��9���.�g]t�&iwy��>?xs�SB&T��8�dt�sbk��Z}���]�-y�|�� ���)Y_vY�gԕèA2D���y}�!z��,���1��8���}�;�w�ug@^ըI�0�����?>���(�i�&�A޿C�o3�Πq�����f ��{9�BSzK��RL`kA��|���޾s��~�j���x�%-��Zz���_�	�������cfG��я��Q��U�����W�@�v !���s�Jpd��&twY�%-�T����������wz�䴶Zm�4�5&�X[[�;H�zG�JQ�9N��.u�#oH�-.��O���EB�:�qA�w0e����N�Q!�,>�H�ٿR;��P8�(��C�R-9E�K�82���n�c��/����_�O��O�͵�}�m�j��=Ϟ>�w�����o�霾�(U�I�p
�n�kn�z�����,ׄv�{Xզv��VD�Eb���yYF��Ω�0�O)JC�Y=��s��>�!e��nVq���|��#g���}����3pe�$!*�E"��-��K���ٔ)UƽbPT.�i�`�ޢʂ��V�٤���R���myO��>�M6�zk4�%�0J����x����$�������� !�R_-P�N���D7ݸ`�f2�V��I�N�T��i����4�*����� U��{��T�uJ�%(�q�k߿��������^W���$+h����9��e��O���t�pt�h|�V�&1	��W3���G�e�t6n��$�¶���D��2�]`�������s���m�ӡ���v�S��q�k
~����*&�	��^n�TV����Q��^�}W���6O!�t��F�h��"o�ź&p]��,gms��7�*��P������Y	*�;�`��>o������Z	�.�8;�уǜ��,\�����ӝ���r��E���������{�E�t2a:�b��V����N��Fb2��n�fkg���-�<��/>��,�9���DY��Zk>��i���W�]�VƬ��,� hu2���mm���esm�^/��G��GF�	T�bQ-�\����ǰ����������y����B'h�%x��ټij��ڤ�A$���N�,	�vމ\HJL3FLp��IIL���Q%"c��Xg��1q&X��K�窕�,ƀ�
������چR�w��MC|��m�}�Ngc���8�ء�f�6�޽���g'����޽��۷����9���<�����,3D��K���@�V*���	�3�qd49�$��qA���yJ��Z�V�6B��|��%'''��q)�h�]���0�8::����1���V*+����{��4Z�$�։�i���A1��c��p�>��? >\������'y]�����n���@��R]�	ޛW����4��5;�oqz�#z�d��6P"�9+���?��?������������z�����3���6!��	���Ңoy �dCp� �<�W�'�����숃�,���2�Q�)����%��S-ב��E�ƍW)�
,�.	v�h4�����l�n7#�r��y��HL����(_�����������׻��j"ˢ9��5}���w��B|��k�RB�bk"�|=.*,sa�HX5�}�E��e(T��������`0��>�$�h�|^0��=�[�tY�3N�^������׿��0�s-�$y��t��W�p����4N��K�B`<q||L9_0�ssw��`��"{�>y���pȳg_������?���xF�b�%(�,���'�s�v�fk�O���LB��1��'hI1�Kj$�Ҿd^�Iۊ�{�p$1^,$i	�|���QQv�iuԊ?i��:��<ĦPC��$���h�)Y��q�uAK�vY`�����Zu�u��^�H�;��c��Z.�%''_<cVN����j�Ij���I�ZX7���ԾB%�nhiH&1�f�p.�DΝw5"	���
.��8|򄃭���5�z=v�n���?"Ks�o޻���-��.�ل�O����CF�<Y�!1�9*a%f��`�!���5\ښ��S,&T�ʥX��ϑ���xo�
噌/9:~��'O8|�yQ�t�h)-��4���j�q�"�R�R�D�\������%�����u�*��	^��D�J�ȮJÖ��y�ˤ����{z���/~��W����?���h<>Ͳl]'��^!��#ڈ��Z�e�Ue)W}KaLs���t���M�r��~��1A+%Ai��!�F��y"a������TR��u͙������IxM�
�L��S���b@y�R��huKUL�O9?;b:�E�B+�HҢ��dk{���\�_4Q4�@�W�I�o0~�1pVJ!A��QU%�٘�x��fT>.5��.�:�+b��9�@Y����7�����Ѷ�Ղ��A}Q�xƇ_��ӫfԣ�Ҝ:D�x��(E����(e�Q:�3X�~���]�I	�Py!1-*;DDa�6MB�縺b:�ɯ������3f��		����_v��I�1QMmd*D�V�E��A)E�=�E���;;[�Y4^���(�Ŕ'�>��ɣ�py�t/��/:`�x(}�����,�2	)�)tPh��i�D�_'�x^N��iQ2��)�%$����c�b�Qe�!(�.T��:�o�77����`Xb@�53�f�Dى�%&r�$P�|(�PTT�)ò��:z����U�s��ZB������ٳ'�������!H�&�A)A)�ҁ@���2~t�6��B䲪&�'���ޡ�4"�D�S#xWq9<�<}��v�[Z�6��?��w��更RE����b��/x��g�'8_�[,:�x/,=���F録X0:�����O�YR��-XrjU������+�j����t���H�I�ީ�z��cV�E]a�IB]�WԐk�kR�^����υ Uei�rc�$A$/-A��}���L�<TU!�^O��n����A���T��dY'�z��ӿ�ȏ�u��%�:S�eVV���9|Ղ���WH�7Mv�
lcB�""��
<����+k��V\��9��#>D�Y\c�-#iUK�7�݈`�EU$�;�lz���s��ȩm�h�!o����e}�����$����z����2���_�o=x�r�p8d:��� cZY�~-�"B�jJ^ݑ}��s�f��`���L��n��x3/�?p̖���j�7:�t���л�T� �HZ5i\�y�j��q$�$	:i��Qdy�v�M���jaV�(�Ap$IF���:PU5*8�/Ny��3~������)�t�Q	�����I�&��x���hcل(Qe"�Iw)��bX�ɑ��W�`H�൥���Gǃ�e<<"O*
���:��FH�xm�����<Ƥey�Ea)m�V��m��*�(�0Z#�B�cr9���/N^2�Ϩ�8*&Մ��2:4�Fŉ!����
���� <4~E�6�RsM�(��@��D�T@+��btq���Ng#��Z���sM+���|�t:���X׎����.�gq�e""�Q�DB�Fi�I&�
:U�<���m�����I@�L�J�&<�q�W�gCN���O;dY4��Z9k[�l-��������/���Ǐ2��"(�ƈ�#^����
���E��<!K�Mk����G����C&�&ic���lؠe	Ҩ��5����(�bm I�>>Ьe��kJ^��*'4������Z��U�A�އ�u��e�
��
��V�8��7?�:yxy�8__�닋Too�rx����;Q�����!�j�8rJ����[�B?�1ʹ�Tu�TUi����s��2h��
��jσ��}���B*Jk��VB�j�oz����^��Õ[� ދ���-[�W�9ML�pED�DS,.99~�'�0��x7�t����8�h��u��J��l���q�4&����i���l��Y�,[tL M���}�,g6/vD�b�ثuݪ�V�D��׵t�ո:6�ZA�#��}�`�J�-V#��AGT��f�7F�e9�Ic"��h>�tT�zE�^%�i�Uѧn��c�(�1:?�����GϢ��GR!z6�i�1�n���5Ƭ·J���ʢ����GO����$o�u7��v�R�Ep5�ٔ��3F���bM�C�9�I��k�$(�N���삗����<!�:EEQV�N(B75>AH��_I��H�x����_~���h�i8<�S|0(�V�N�G��f:)�6�/�ll��1㎈���(Y��b���hţ���|��ƀ��aK��hƳ�S>z�%�ш�l�B˽�C�A\U�r�{�L&��c:u�%��(<u��h�:�IS�iP~H[1%o{��x[�G�(ݼ���K�; ʡ�`�soy���wYT���$�:�
X�N��t���S��O�m��$��x����@�%�ɬ�U[�<#1m���*t+mI�
	<8���_c&�u�B�����l�٘]�VYnڜ�]կ.�W��oF����~��)x��DEDi�m0�����|��ϊb2�v����)��]z
���� ����4�x<֭��ot�_b+%::ŖE��L��^�#�-���"�z�[���h���XV�l�F�Ң�(Z���������^��+ct��]�Ba��-�4I�}�%M<��-0J�U��&��{F8Y��JS��M�6�������./��!�$��ɑƻ,6A��Ҟ�.���C��Nא�ڬ�Ek��0�̿
��~�k�f_�����ﵓ�G�xdV{s���+�/���j�_q��o�b�4#����)�ݖjN�5&��Яb-�ق�dĢ���5��k������������UE1��'��Z��ʤ�������fιՃX)MՂ�d���3�=����q9��]ۤ�
k���HM 5B�
�!k����`�ńZ"oL�mZ������
cbsrt���G̋���'B��D�^C#
%��L8*.�#�ʣ��Y���xhe	��wnߣ\�9>z���|5&�bJP0���L���a\�XB��傋�S��Oh�����o�L�V{�2�sqq��:��@ek���.P���
-�o�˫H���1'8�b�b�=`k{���]���i��Q����7�X,JNG�J�5�]�������z�x�s�P3��<;z���ǤiJ���h�jŕ����%�|F���q{�F8��F�6F�b��b����t�$�ps���t}.//լ&���;�6�t<f2�dQ�i���-���=K�]fl+uM��$�HC�_�ZYZ.5�_���⻖������	��|���S�|��I��Å�^�?6J��'������f#�pz�~���?��������1���E9wO�q�*+ŢJ�"��f�?���V����^9Y_�u7�Ʒ�9PJ��*4���('���̿���^/��T$	�DB��κ?jIY����Z�W$H��ؼ)#TuE1��=�����z��\#��m�����B�eE$�/я@l�L"�V#���Y�I�����A��g|6�[�v_�.���\��;-2�F�\�7�^V�+���b���D�E�Z,V��Չ�ʸ+�4&�:o�����(�'g'<{���'���1I���6n����{�9I kKL�$&gmm���5���UAY.�E� 6�������r�~}��\�x4���!���>���#�<IQy��;�c�bVVܹu�!K2Zy���Lo����EM�
�3L�ct�w��t�W�,�X__����z���K\ KeI��rV���x����.��%Y�C�d*!x(��ɘb:a1_���Nw���w)���Ֆ�\D�OPH0� ѓ0�wK�P�ӨA�;|1'(�r���/��i�LF������~�ڠ�˗9���6 UUD��tJY,"�aqδ���B+R�!h�7qC����&a���`�?���w�����bm}��o���t(?{@�X0����b��2"�w�v兠^�<�����no���Gy��f��<}�gϞqzz�W+iL��xo���q5*Tԕ0�sv|D'KI�gm�����n��[��ՆO�Q	Jiʲ���'O�����OYT��}�Fk� ��gt�ED_�&����B��Y2z_��yK�Jϑ�D�jU�E)��4�`���Y��cv,�0׋4mϒ3��(Z�V�_tC��{�%�On'm��u���d���Jkkq��lj�Z�(^�̷��~�K�~NW�h_�zq)Q!���Q*�J�|��߿/�����>��C�I](iϕR����ת�-�j!J"�D�х�
ثrt������j���>�B������^��;o��BQY��6��������S�D���$11!�l�Ѝ���c]�u���
7&��h�������6�OO(��t5޽�9Tl,E�>ٲ���ż&�ID�p�nB]�e�FQ7�Ө��RW.B�ί�4�4���\g�'-kG߾łn�����[c2�EkMh�8�[!r�.U`y;糇���������i4���<~��gsn�Ϩ����M�Y���N��O~�3����#·�r��Rʪ��KT�"�߾��![�&f��g�����j���)UU�����������W�LQ:�פY�|1���2^�xy�_Wܺy�V�!o��w~��`���]l��	E�qV��Z^�8���%7����	���m����4>��cF���b<�ɵCD�%Q!�g>�1�Ϩ���ʨm���ʒIF��|��G�����"�Ak���]�Ii�Z�L��s�kOYG��[$IF�g-�
WVL�#./ǔ��	�����c:t;�l��i%}���u�w眃��eI1�9�g5u]3���8���ϟqyYPۈ�4A����
��߿�_������{j��1�� ��ǻ��=�{���7�կ~�d2i���,��6E���,퉪x�7�[G�Փ'O��w�~7��2�jA����?��������@�c��JҨ�vok���G_|�txNU��[?�����N�v7G�h���Z%X�wn����V���c �G���ʹ�Y[�S�\m)˒�dL&��ycU��i9Y5����7ڱ\kJD�r�p8H҄�*�i��I˪hk�Z���5�����>�&�����Lc��A-���i��m�~�ӟw������mv���o���m�H-BR,����$�$"�����<ֹ�O�r��r�B4�.�Y�IL��:��H�D��!��K�����A��������㏿w�(��z��������T.B�^��JI���?�u��fÑ�*�X��=k|�[TH��cU���/�NRҴ�Z��HCr��6�*ߠ�}�_I�Ccyʲ1�C�q_�7�k-��R�S�Yކ�xl�ڴ�4o�e-"v��[]Z�i�am�1M$MS�xW��BՃ�B�f��|�d:b23�M(�cQ�S&�F�3��9�op��>�kk�SC��S�9�]0�g\��P�|�Jd��e�z�*5�?G�j<:���R[����{��6F<�d�~+gmm�v�cm@K�����zLU9jU1�8=>�r�&��6F)��6*l��[���	'g'���,���"�2�&�b2����K����F�}7v;J���3��x���G_0�[���u�t6i�Z�:]n޼I]͗S���#ht-w*q�y(�)Ǉ��򋇼8���<�W�e���×t�5�Ulml��{��ݽRH���*`m��5E1g6��P��Fc�HL	���J`�����wx덷�ٹ� I ��*xt����l@Q�x�����1�$|��M�5/����?3C�    IDAT|Nϼ,�ᐧO���ssg�b>���Grޠ|W��cL��Fm⫨.����kz����~/GT�(A��zO�bڈ�)�^�;N���H���+[��<*(���Ղ�t�h8$	�Ʉ�(V����=4��_�{�[}�9ޞ�m�(z�H�E�:WՠL��R�?-�������ԡ���N�]�>F���_\Cr���W�ͺ��I�2���j�V�.�^��)�t>����|Y�}=��g�sN���!��c��ޙN�-����Q�V�7�L$s�
�t$!.N7��*s�ܽ:�kIĂ�Z��o�# ����j]W3��V��@i�E�м�u�Ĳ�[�dF���I�������[��{Z5�ߡ\"��g.���G����vz��t:=�2XOK�u�.��-0]p92�Wxp!�s���F���h�2��m��(3\]���Qc뀳0�O(&c��PԴ����f���O���NY�������PB���},����$^�Sj��[��hmQ8_���Y�!��;�yA�:X�F�w�X����[@r��X�̊9��/.y��1k�d�a{��w3L����6;��<9|F���5���V��D4x6���S~�ϖ��W�	*$�ה��U��&��D��cs�M;���ln�@�a�\|�/G�"8-�U��P-x<�3�L8�Q5�ʨl��r�cP�������Q{{�dgR7�  8D*���m��6�8����J�A��"��i]�L��)�����;�i����zl7mJI�C�Ao�v��{�#%(cb���jWOh�J������|N��{����?��'0	�c����L"��9�&x��������g|�EME�7����u�t�,n]���b��H���999c8���
.
��5���������+馚Ǐs9R�q�-J}M+4^�&�Z!P�:ˀs%!h���u%J%�uκP�Y�1E�MI����i˟�I=i-.��M��+���?��%�������� -R�VR�O*�[��&I0FW�z]����t��u܈E:�%Ѳ)�_˧��oЬx���9P[+�7����%"�ޫ���߿>��ÿ���[��W���E!�Vˇ��b��I{���X��~�<���k-�%��ɞA��h�8tX����$�J0є��W��#������o���1�
)�}u�DZ7���t^7On�Zln�q��>w�q�{��khӂԢ�܂��\pt��O�����c���]��ǋF���$�	��5�h���e�b4$ʠ�`E�XB5c|�ç�v�`n�ڦ�O�m�r�U��x����!����.OrdYz���{�="2	$�B�����j>�j(3Y%�43iQZHF3��h-�?@f�ϖ�^i%�dM�E�#gĚ~Uw=�F&����p����u�G"�LTݨ�<f�gDFzxx�����|�;8'�Z��y��:�+:���@Dh����.��k"�8�()5�Fxx�KJQ�F��-n�{��[(F��o]��u< �Y��Φܻw���h@�{k.R9a0\gta��I��̳u�*o]����y�i.)K���+b�kc:K�-�R
���p�.E��2k��oq���
�A�\p$.WxӷcK��V\�T%��P�%B64vE�,m��'O1�[��1��1���[����1���ѣ) 8�S�x��)�qC�b��� ii���*�f;����vΚ��T�6�͘��5����_��3��w>�l(�X4�o�\K�r�d�	 N"F[�i���	�4���G����翡��	��5�!�c���QV{�RX	4��wwB�3&�k�qy��!%�@�az8�����i޿˝�>��'�ۨ�
Vrߑf�!���/�~|��Qvw�u~�)W�΋7�n��@]f���y�����2x/�HmLM(lBJo��?j��vY5>5F+�ݵ����O�d�>�� >�����O���G:�����b���+�;�Ժ�lTIM3[�����d��nE��ub!ʏ�Ʌ��҅1�X�R��K�����U����fę@߭���(�h�h��4�XPe���x_�j�[��v	����:hD�JT$!��p.d]�vI�>��ٿ*3�9��e��-�MSVD�$��������2�_ЍkG�
���tU�!d�6�r�*7?��?���~��K��k����^�����m��u��K�؟Ly�7f'9M���p���:��m�>��|;����fF�5��A�jIi��<݆_H��#޻u��Kk�oq��m.]��<��g���K��|��[�M�Svww���c<x���>I��o�BR�U�%�{;�'f��{4�6��������}b�`�$ib|���/͔0�0���֥.\X�	��X���amT��ŷ-�ㆺ�D1�u8[`m�e���0Fi��w�&�;�Ƿ��w�z�2��̩z'�2�qX!j������u���N�o����SNժ�t̠OS<!Lr���{̏��b�!�������*�������|��`>*>v��C��Aei�	�}�k'�lm] Ě�3��g�lS0*���'��<�������,")֮��F�O�9/A�$�~q����}�t����Z�!�-P�`M�B,��<%E4`D�.���1�����1���s�chĄzU��[bPJ��g:�#�Y��I$��ɴ��G�-�l���s������b�S8���Ң�������=Lw��1�oo��n(Ӭ�O�̧G%b�!�j�8Ve]Y#�u5�����4|�-��?�O?���~?����Xo�������9��5��4�se��PO&��'O6�ww�tC�EI����en�u.��E�6`�qh����%�
"b:џ��T�L�1���/������k:5��ƙ@_Bw��H�B��=]~�E����Ӹ�J1�!�V��Iٜ؂+��&EUs�*LgP,���с=Y������������X�SY}��M�:�[����h4����|��G|����z��%$�Qm�M�ea�8b:�Y�ؤ�z���p0�&�U�������Y]���O��6��^��2@�1��#M��$0�3����8�Nx��7ih�7��i�u�8k�i���Jz��m[f�>�W��'������石��Z �^S��)O܉�H�	��=�ٲ�����C�Z&��G�~�d�MJ�%I�D-��{�l:�`o��G��y�W�^Ŕ�<`�����ȓ�S.]�`4rԓ=?���_���~y[s�-�C�%�W�t��<3��9��������;��F%X����Z+m}H���N����.��?$�DU��5��
�;<ԓ�GgL�O�N']Ex���͔�B�ޙDY8o��`o'�EM�F��)����������{��x���6�g�4�Y�+^�Au�?�X�f:�Bw~����Ε,*��\5�ӻ�.c ��ͨ�MTeA�a�k3[ �n�h1��jn��'h�H�"m8Z��s0> ��ԶB4g&��ۯ��x�YM���qHS7<Y�I����b����|��|̅��
/�=+z�X7�	��x��g^�+��j��j��N�)B�FA���$�B�	�������8Wa� }��'|��O_A��W|�O������'�Z;M��ǅ�ֶ�ș�Z[��¬��{{����Ҷ-�ᐶ^tԀ�E2��dڏu���L)�jV�cz.Ѫ�aT.����򓟸�
�oO��FkL/������Ǒ�2a��K�U�K~~�ӑ�ib��e��{�M�����E�tMy�:��X��I˞ږ���o��	>}9@QW� tm���Cd\O�I����0EC��)���eg�)��Ɏ�H��~�ij?~̯~�+�<���o���ϙ�p�|���"b�1B
D��:�������<�~cZv������LC�s�ٳ�,9���f�����p������MӐb���t�Q�&�B�S�*�����=�pv�W�Q&��_��S��Tw]�[���L����s��}.l^"Y�`<e<��g}�2kÒ����gw�.O��gz�K�BU�C!�x(�l;�}�8RPB���f��?�*�)�1������|����~���� _?%�O�O���Q�@�DA\�X!Ɩz6CS��䰻�)6� :E�DDsG�f8c(J�T�^hSM2UK݌��W��!�m���o)6�EI]7�Pж��aN���C��RN���C��b��ռ�p��f#]�UL!��8����:5�K�gP�XbP�5X1(	M>��IH*X7@����b�Q$Ke�0����̅����-޷�~9g�j����]�[�����O���c����is1/��: 5�b�y�W���fw����[�1ѵ6�V�vXɪ��Ŀ[8[��u2����a8����G?����_���'vs�q��?Y�5����?qI�'�A1����4m9>8ܘL&.�,�D@��<�I��Y���`�8�f�����#�N��T%�:��lc*���*$����3���s�U	A��$Uc�(�|��E'�~��S����C6t�Wg.����8�V)�k(V�#���2�޿��8�qٖ��U���~���k��o<��_���t��*�k���f�	|M�cB}H�v�<��d<g�g988 FK1(1����;��1���~������|����6t�-��Ɩ'O�p0>���#O[�3���-W`��6�:�_7��V����>١r�������JLk:��k#�@��hB�p�ϸ�	dm`)�!Ea�}"�-e�!J[�����c\�&ԖH��!Q�1��Q�QڀȄ䧐��I!���1Xk��@���)`�Hg:]O�k���r�)�Hf�А��Y���2�m��bPr��JT!h�$���qW!D�`�v�#崣��H��F���lJHu��i�mZ�R�1B�&Q�HDf��WLYfB�<�u�o�o�{q���,@U�o���b����͆�JW@�L�����lC��l�}�I��M1`�ҕG*�mC@	����{9�|>F��F�9��YK���/:0I�d޶-V���H1��L�;|\��*^���>�;vrn�[D��Q/�$Ĵ�
{�IBJ~�!�XSUv�&L��OJ�X����~b~�㟙���gG�1������V:w�R�ܞ��c���z�Q U���Q�g͠���Y��#y1*2\��qQ�x�X�Or����j�uSծ�KlLq���`/�n���x��,�O�����L�V�q�&��5	�N�-�XTɓ�Ƣ�U$w��<,�Эf��)�m����Z�F��lfk
<-�Xc+�t<�Z�����%�P��w	�RT�v���e���>`K
r�1M>8�*�4�1�3p��{�7f�ʈd*� 53��Sf������}�n����1J���8��!�<��~���se�*1���ȣf�)I)�6?15����ȕ�
�1ⳬ����;�[��bp��J�9Mn�RPtm':i�j��-.�rv>y^U���sʪB"[uV�i�c��l>/H!Rh��~�ՙD$c��su\�P���s�6B؁�C�����>R~}вh��#��0L'm78J�Ďc�1� ��@Y�m�����'H.͏_ �ݙ���EJ����`�J����:��^��t�-�o�!Q0���S����k�':�N׵/1�<g�.���UC*����I�4�'����˔U�82��{D��k�Gl($�^#��WgX�Ou��EP
F4��巏�Pu��q.%%H�R�5�[�H����I6W E�y���\���������7)X�)�|DT�K�f�W�RJk�&R��f���؋&��0���J[��+��O�n�?�ѧf��j�w�����S4w���n���'���R��*�K�1�}%�������U����d�1�r������A�ˆ�>t��������?�Ʈ~iI=Vk1)��)ϯ��Q��L��11)��@���Jj�0Ŗ�%v������gc��U:F�0&%!�u1�d����u�?Z��7�JB��}CU�y���(�������EvN�/?�wqH)Q75�{{f��q�����n�V�����
!t��ɼ[ċb�ZK+������r�끗�*(�"��B�٪Fcw� gW����i�$���V��G���O��8�~��U��*Q�:H�Y�;c�F�����Kg�.�5��O�wf���p��7>�[Ě�K׸������>������I���6�E��m��(T��!������]Cz�0v�XhQUuRu�Y[M7�f6�!�)��d.��^/Y�u������t���y��������^}ߢ8[!�z�=
'�ݚD��d���_�+8�]��Z�I	��]X�8�w�����S�5M�d� ̭WV,Z,I�-W�j��X��+2@��<~����]BH81E�1j��@����!/^dss�A���0�����$3Σ`����O�ǐ-d�h:��B3k��$�:*5��XYM���2�8
0^%�8�����*��i:���y�&��͓�����1W8ۈ��v���%�d�q��GEQ�����ч����_�6������U����pq:������z�O,l<']��'��>dk�謽��dR��ު�쟪�7+����!��)�Z�j�4�l4�N7Ƈ�E�4Y*�V���ŽesW,��E$��I�(DT�ALix���'v^��-�3rlI�HL;/�:s,"9����]��RM�QJY���֗���A��>�X�*@c-�a�h4��+���kvvv8<<̀�Ȃ���t��]ڼ��o��[W/�6Ќ's�O��B_|.�Vy�� ��++)!��*�3�v��\�����A�eA�:(8��������5����?����o��=��~˯;��N0�����4�+��ê*�Y�F�U�O�[8�/[�M�?+Fͧi���TվrՌ~��?��ʁ���w����?���>*q���?�,������U�+_i�FwyjL3S����b+�?J��7��w<�[냑Sgdm0l�1ƇP6���Y]�O��y�^�ڟ�Si�_Ac3Ţi^@�C$��%q8+��ί6���<^y�Iӷ���$�I&�K"&i�����`��;͕&b�nA��� ��a}m@QX��Q9�og��<a{{�}���x)2UE����K��" (Y���>�r���'�������VX �$Yk��9�|ik��׮r�������Ã��2O�+����N��F�����lQ#�pe��>-���E!ar��ף�>�W˓�d�NJ/����4�uX>!�k�$�F�Q��j0��?��sM�j ��i�Q.���p�P����Ц;X�����׳bˇR�n����z�%���vZb\�&4��8w����}W�vW�ߨ��ٌ4���������
6S9*�5�~���v�b�Δ�rMqV\ҤҴͰ���tR�,S�[u���h���~��@5%$t ��@Hڦ�T��^��|����:rxo�Pp	�6%HJ�uH�9ӷ�^~*ɵ�BF0�!"�͌���\���/_b8(�~��Ç�~��z4����6j}��%�b�K������ds�kX'�f-��v��E��5��iU��$B����pĥU��qx����cU�'��42��v���i裐��T����x��_�3�|���q����*Nf�~w��� �o&�������災��qϩ*Ei��i"EQu�z�m�Uj�Z_ۜj�֕E+FRR5)�.!}��	�}��~
��Y��^/�֤Cm�P��G�!<����ڎ��ҍ�{ab�nĢ�k6��B5ҡ	0�n��6v͖���?֔>H�ه�UAGU5�UY�\TM�o�Q;�mx�}�ڦi�v\���(���&^������R�c�6DB�F�[��y�o_�	�ŵ$d+�؈:U5"G�ď퍗{���;��#����"]C��K|��;���[\��"����Gܿw����K��}ȕq1k�b��(��P5(��Xc}4��'���=e�`/[6��y{�{*ٹ�ϻ ��    IDATH��Z�%���鄃�]���2�N�L�T�����Aa��i�Y�TL6}�k��1��'ѐ�0Y�>\���4}��e:���E �U|���y�5^���_�G�"��Ѣ��N�X��DFeYVj��� )�PT�ںn�1�^5����$�=I�`�Rnc���ZQ�E����jU�q:L��D�Vn�GFt+Z�D��tr	�+Q규wkɷ�c���n8W���Z] �@<���:F?�L��I����t:z��|�nKO����{��.lI���FB�4��U�I��1\��~��� �-��i��(`�}�$�dR�6�/T8Q�Ē<��1	���)Pcx��5޻}�wo\g4������#�>}�o)��ި�8�̲)����F��P��������YSO���:#Y��-��N0I��b%kg(��Id��4������H52'}+i�#^ F�bD���J�W�e3ꤽ�����w��v_���y�&��b�{�%215�Y@U(܀�pHJ	��_��E��u���5]S����R�B1�)�!�Ԋ�Z7j̄H� �u4^ ���v]�#����)m�&�a��� �c5O.���cw��/��2��\��-��\���E�����B!M�b�{�F�|��?8g��MqЗ�>.�X^�d6E�PD�pe]W N_��wOP�ڳ��FM�2\[����*�!�W�)x��w������7x��U���޽�l?~ȓ�;��I$�eF,���	[qEE�F4m�(,�{�ׯ18,���|��_�gUU1�L(\E�b!��RG�+��	�ʕ+8������W0�1�\~�׃,�
  ���������r��Q�ٓ�2 㤮"�������<�D�wg�A�	���q����}6�s{���,Kʮ7o۶�I�vZ���/�����糂ھ���kW�ɯ4��L심YN)冚��Wg���.8"٨:!�h�����{ՠ2h�j*�"8gP�2�Xi�/$R���V�zM�Ψ �
�*;�ͫ�%O�����P8�jJ���0�8��l4kf.���s���ׇ������;�eM{	UW���}v�(�K�l&�>��\>)�}0���ӟ&�����[gb�Jk5U���%f	��Iz�>�~�㪪HbH�-iC.�غ|���y�;�x��UF�����}u�P�5�]�_�N��j�blژH�FL�ŋ�q�m޽q�A阌�9�ߧm�DB��ш+���u�(�BdPX��u6FCJ� �L'�L�����1Z��	�t���fiۅ,�Wo��t�LC߲k828<<<����8�}.sx�at1$r�a5��<��E�)x�Z�h��(E�*I��S����El0֥���8��AEDEcD�dj��q��)]D-�4u�&��!�!�*xoC�4�r�Ƌ�u�S�����Q�1j�Qb�x�cw�)��MN^���`�ٲ��ֺR���}A���XN�������!t�Ƹ\�Q�z�&|�޹q���!m[s��W|��_���}f���a�D���*�������n��wo��kW0ֳ�󘇏�3����1FhB^iI���GX_��z�*�/_f}mH�3&��1��H)��p��/��=8�Mq�r��z�
����8~9zV�(���k:�3�Fͼ���~ Ů7�t�|�ShE0�řO��[�5bR�)*�@JEU4�I�Ģ�k�.�;n?+��EPє��dU�A0�{������p�{s��߿��Y?rQe�;���\��N�<ޘ8�{\�+���M!/uu'����5Ε`
\5��[7���l]y��2LǇܻ�_���ܹ�%��!)eX���	\��� SW�+��pĻ�����=�~������{<����l�%kQ��I�jD�ź���$�j�ƥ�Wٺt�����a:�g6��O����g�!���P2�v�v�V�|��Y��x��h5e�c	�'�E�ӋS���X>7G��]�����}�CU�G�f�y�Ҩq��������+FZ�5	�$�FAS���hcD-�I��,7�l2(J��������rG�|���ӂ�ש��x���`�1�<C���!�կ����gf����RKnM�]A�Iz���j��h�(�؂ \X����~�ÿɥ�ˠOy�����_����<y�M���j:���C����9�5��ܾ͋�����ryk��-���<|����'���]���U@=V�`�)sJ��`\6v����>�Oi�Iw#�\XqV���g��i]l�	����c�oE,�{��ih�����ى�П�k��+�����-ֆ���;Q)�B94�1�5�1-��`:�*kr_�Ō�<�Dke��]���5�B�V{����^���sm���?�J�"��:1�
�&����˷4���5��j"�eT2(S<]�]P�P)%bR\Yq��M��}��Zcw��|��o��/Ν;w2���PK7X/��ՕZ
g��իW�y�&W�^�,�z����~�ٴ��˒f1|���N1�`��Rĕ��FC������d�����b<U��G��J�JZOڞ��{�}ľ��w��}�D�D���g.����)�+ˍ?��`��YW~�Z�1�3,)ET��Z;�Є�[P��<.�`qe,�Cմ� ����~r��<�e��ke�Ln�YΔeiLW�e�I"�ꕽ�y|��L9�*
ߚ^4yU#�X�dR����EE��X���L&5o��ۿ�����Ν/i��c�
��v���T��\�����n�s��tL&���=�7��>�i
k�{h�%F%���Մ�܈��%�]�εk�p�Ѷ-�Ovx�����pn�g}	Ë�Az��㟷�J*I����������W���X��	�������%D�Y���[��3K�v���8A4�l.߿��x_�C π���U�a�x���}Z�3���{��&vټ�M����9 ��+\��a��j�M����� �㍎3��Y�)C���J�b$:�Ϟ�c�cK(˒<@�d2k�������9�?`4d����5�Ic�����[ܺu��W�������Gܹs��;Oh��Ҭe[c(�2�#�V��x�"��~�o_�(
�Y��M�Ǵ~�R!� A^A�9���j�3}ov8����=��nguss,����e�y�=�Nd?�U�K_%{�u���=���m����Z���.���4����z�ε�0Z�I�}ǹ�,�g>��8F���8W`l�ֈ�5�	��@��_�}�'���8��#$I�Ĩ��Q�ѨI��6a)vb��� u�>��B_i+ �S���&�<^��?=���m��wvA�J*¬��D�x������O̚@U��쀠`�a�q��[ܺ�[�(�I�<����|�)���S���`��QC�<X�X���Q)����*�X_�k�����/�՝<�W�]E�Y���t���a՟�ϼͫa��������S+��x8I3 s�`ur6s.u�������wr��<.��f���7�_s���v��'E�w�y��O!=+������7�#�d��ǴB_���cN2��O��%F�U���ZO�~������IX�-tL�v�M���Ο��Y��;�,�Wڑc=p�}��N<[��2>q'�I H�\?��7��z�K��)��x�^�[#��-6�礟S�T}V���f�g�2���Y�>�E�j��"�=�G�`>/�Zͯ����[f,!�ު�tm}��f��pΥ)����v�j��ε
ߢ����'PL���|���*�����}>|ȝ;w�]��SU�gQ+F��p=�L�ommq������u�666�L&|��W���?�w[!���tt� 1yF�7o���ߦ�*���r��]?~L]��f�\�����߆X�p�N���~�-H��y��=��޾�����ZyrtBx,�|F%���O��߅.^��~���=��n�>���Ua����[|�c��҆E�/��U����M��,�_g^�Ǖ��� �ˎ_�;�qΉsN�u��uZ�����������[_����O��G�7-F�VEE� ��r	�Y�}JJX^]�̩�+����}�n��'hBU��!e9�m2X[[���?�>|�ׯ_�ãG������/x��q���ɫ��Bm�^�o0�aL�h��͛7y��ﰹ��d2a{{��>������4�{�@U��6�"s�on���e���Y�d����X�L~�3kF{;������߱[��a�Dt��Iz��d����㣽��n҂e�N�!��g[�*�}��l���&A@���nU㉠�E�A���Y>Þ/�c�AO���~�o�?�	�y��q�Ӥb��eP'K��J�w��V����cL""�\a��1Xg���f�{.���;��g��ŵ<�%��Ր�GE����VTU5_i�1���
�f�F��v����8\�(�� ����&����G��7or��E��}>��s~��_�t{c�����$h�%З'����Wʲ��[����y��m6/l�t���`�����Oa��sߞ3}G��ۣ�^g9r���:�*�B��(_o������:H�Dn�t\ ��|�G�:"$zI�2"�������j&e��벤g��N���.tvϜ�%����2sܛY��+ow��'�Ó~}�ذ��>I>Б���2��S�����e_G,�w1;h�􄉱��9S:�ֈ�^ӌ���'�g?��Y���7(��������kn�E?�b"V���?���aޝ�B�Az��:?I�H�m�1�N�!�u�oB���o������;����ŋ�D?~ȧ�����/�~�F�*���ӗ�ж3���ck�"7n�`mm�m۲���xrH-�r�u��r츕ٷ-���8��g�o��W��93��m�Ukw,_kk^��<y�Ư׳��������g{����ѕ���u/<�f̋�N��%3��9�*��%��J���LO��=��;���<����q,�i�(���Eq��x����z��獛}���U+�Vމ�Κ5��5�����1gouߠ8[�ݢH	lJ�`,�d��|c)g�5�{�s8W�W�ٳσ�&3��^}���dp8��p.�ԂZ�p��%nݺŇ~ȕ+[���y��W_|ɝ/����!�� �ퟮs��|��������?��}�֥M���p�����rZ��x���m��M���c������� �\����X���z��"�x��BT>?h��$w�:��L�gX�W�<���3�)�F3S*Bf�̢�d���*�3�ǧ�O�J>(DMWh����J�m5�������~��p�5�Gu\���ī`�����^��ιcu½��/ɋN�2~��3}=��3} )%��.2�IuՕ�!�J_���/�E�g�g��
<�oz�	���|�.�n]c�4��5������@�����v,�8.���F�2/�7�t���\��1��Xm����p8dww��0�����f|����E~����e4z����~��U�i;cP�q��{\ڼ��H�6̚)��!�������]�dQ��%z֖ q\��i�h!�|��&n��8��K�z���>ޕ8���h�:�x��ǂ�[-�XT�0��^?�>��`�?~!(Q��,���*^���4��o�xn�����vL�1�9��@&溾�LW���@/<���7��5͋Ɏ�� p�ƋX��|?�}��3��2�{��nk��lB��Ĉ1QL(4�ʵ�����y��ę@�A�ɉU�D��"�d^�:)y�������u����z�*�������s�c]�]��bTK"֔T�u�p8��W��x�ob��`Pq��%޺z��]�^7��)�lK)�A��U��>�����_��_��w��`�x����';s��=�r���f?��f��:)��0b���q���Y��*qV& =�͸�N�xFW��
0����XT0ϋ����Ed�0'k��V6јȋ
5�=��~�Ȍkϼ��~��ǅ��9��90[a:�/�u;�wʉ�(����۷E�`0�,K'���Vq�)��y|�����q�����q��Ό�`�w7�ɈD1N[�$C`��r���{�3��ٺVZ��aJi�.���b4�{����2��_��'�bLs˓����yY�x��������ܾ}�����r��=�nr�)��*��[J4	Q!E!%�A�d˖6,,)$��|N�>W�Un�|(s5�&8����o�q�-�~���i3f����Y�|��OO�SwmI��~��
,L�v,*b�-r{&���������q����o�3��ߥ���TP�2�ޓ�Q̯�����:4�4E���}�]Q�l�_N8=/b5D�6ʲ�G)�:k��Y_��o[�FՀ�t�`�(
�4�(*Tc>>���!$R
�k��q����٬�mg��e*Wa
�GЀE���!N�X"�f�w�p8�mj��2�͘M'�豦�үB҅!oǀ�����%y��My��!׮]����?����u=/2��)%B�\K/g�?N�������|G�r�`+��:NwgN�W�uW��>�s���x߫�a�x�[. 9��{�Ngh�c�e�|!�е��DD�X+)E�օpoc��9%�-��i�fE�d���f)�&�Z�^D�r��Z���d�����۷y��	?����������"�7BϞ�Ч�\'@�H�!��	I��l�Rpue��?�ՔMl$�ّdH�`PJC���q��gO�9��#Ƙ���G��ٌ�F��⌥��X�4&�&R���!	�*�2�̍�B@K��A%a�+[QC�<p
T�+�d�`l�MCUX���/Ė���p��0&���P�:B:�.6_��A�#�,_(܀�j���W.1(]�ڰ����A�A�.P*)�"��#	V�,q�0k[|��x����d����F����t�C��p�2><d��C=~�ݯ�dg{�Է�R!�|��m|���{�_�N&=z4����<�GZ��k��}��܆�cY��鋗^^.k{����}�_�g
U�I�y���)�0)xx��b�ř@_;D��+*��;�a^b��%-m�.tƂu­���C�Ww�`{�EQ�������Kz�QG���&�������RV�M��W�^��$_Z�,n�UJߚRW������ɘ��`I+=<�������>m,�����6`lg���5�ѐ���J:�)�Õ�XT@c"��E�G�쀌���8ہD7}$�u1�� ���	!q��8�`I�����pPRV����䐃�]��'��|2�F�g�k��$��Z�ZT#I-��z�mnݾ��k7ؼ����pP�֕���iIE��4�.��*)F��Ě�l�C �@���T�ӥEQ ���T�m���Y=�+L�Ϧ�v�{�����d�`�z��2�t���O�}o_�������m�+,q?n�)��q�8
��_)��#����8fO櫲���{��y��V阽��E�ͳSG?��N1%IIŘ�ˈ��%�ŤP�&��s��-��߆�Od�׿;
�fC�j�>���8z#/?�t���{�q��E�������]����={�c��j5PUU�t���3�58�0z=N��L���oy�fm.�*������{�r]�4j�V��|ٳ~�q��I7hb0�@�E�ePٺ|�w�y�˗/�\���81����`'S8J�8�N��� &#*W`
Ga,�C��R�v�
+�Pƹ�bĊ �RXK+Î�2�W��1=ܣ�M��_�����3�ݽK�	c!)�W2鉭>������r��������K[����&
+�X'x���dM砪OU/�[[�����l>ى0�-X����Sȩ�r�ƈ��d��c���K&�CrEr���ު/�s㸔~ߝ'��q�ެ}����.zP�0��;��X�[8��yR�g��C�`(�b�Y�:����~	��Ԉ"��1u���Ι��<�aq&���j�J2h���Y���S�g���C�����6k������K���� �� �o�DoΜ+��Nu�    IDAT�~b�t��-ȀO��u�EG�gW뫃Mh b���ƐR�Z?C̳��E����:�~�cy5�� Y# �5�߼�����������¹��Y��0�m��ӿL�SЅ�����K;k�5�����93h�d=!BH�	p�r����e!(-)��+���3(+�z����������}m�C�؁"A�d0����[|������w�JH��{8��$c;p'���c{V=����wk��T!%Hm���&��,WR^�AE]�L��y�����$i�$�C�D9�����f����n�Xb�z x2pXf񀕖��鷾S�r���o~�����х²Fo����Ξ����>�{��)�Ŭ��󽐀F���ak��oz�q&��xo̚؂�u����E���X˫�eEJ���ڵklooc���*��)�锭�-��X�#�1��~�%!�Y0��������7e.� �~G!���I��D�8︐o�g�=]��9��2�e�Rg�c$a�8Z�;�}��?��ܼ�n7��-��&�0����w��$���~k���|Uf��ɶ�vђ@�#��2<7m5�� �QNhX ������dXMK�\�$�Q�U���s�#{������dVeuߪY�d�s�9'N���X�[���8KflB�C���`|~��?�c`D�T��1h��D��=](BU�)(	�u�%t*΂�w��!?��S�%�m�	�)�yۥګ��H�J�Đ�3�pr�>�l���ږu۰Y]��\a����)gGt];�],}uCUUx�ǂ��9�v�ۢ>�FXT3�K�,��ߴ�]~�fu���
���r�{��sr�.��,�Ec�Z?��9;A�D�u�İo�>j7E�4}��4# ���_�M��LGz���ϟ��y��@��T�=�g���@	U�mۑF0 ��V�?_��-h.3c7WWw����V����f٭z������3�EU�AS�2H�w���)��r��M��?���DY����/�3�2��j��A�&T���ВĚ�B?p�y�ܸD�0ҧ��$���B��Z��ڍ�����Ik,V�3]�wb4U6��ng��{c<<�*j���ܽ�wN��\A"���-�͆�=.�(�|��E�DM��.Z��'��ɳb�(xLヨg隖���eg�m�����ق��i�5!�d.2�g,Y�ʲ�,K�ީq81D��V�k�t<���6�e��X� i~Eeuu�'?�	?��_��ZQ��|�l��ݎ�n����iƍ�9��n���u��U��m�^������Ȭ��v�_^�ێ�m *�|ƃ{�y��#���������yA�X��HBL�(ߐ�t��~}�����4U6�߾����noo���2ӻS�~�y�c��(�1��nԑ�78���c�}�ѽŶ֎Ǹ�M��a-�1Fڪ�1�M|��wX��"�ҧm�g��ɒ����cdou��m�VUE�e4MCUU��.(˒�(���O�{�xæ�{���E��l0i;���'nR�7'�(�L��5�C&tB7��!!�q��Ǩʻ}ᛲkW��*�O�Ӭ��eYZP#�UΫ/y��%O�>e�^�c�\2����}H�գm{�lY����� �����v;b�cZ��:��I�SeWoi�5yn������?�Xi|U�!&�k���"�6�>R����(m�u���:ʲ�w��}��������3�2�*s\~��n7��*�2�����2qз��Ib��뢌,yq��8kH�����sN~�GGG\�ڂ��W��w> ���/��/~jbS�g�T�s(0�w����c���&�L	y�����l6c6���y�!�}�@fzb��X?$|� �Z�EQppp���"���%��_�6Қ�y����V�������l��e��l	a�FC�T25Q1� VL�$�F�l�/`��-�G�)��]��0��-�ŌˋWj2�db��M为��u�!�	��O�tp*�Hw}9�n���L�J�l�ح5�e�Պ�jQ	]�fĘ�֊�%=��a�!xBƔ��"D��;����m}�)&:����Q0�Md�k���#\�!MS�n9\츸�S������_��/{��"��Ξ�}�����ꞣ���@`l>0q��آm��)�G�T���l6�N
\~���.}tD��8>��3���M���"˩��3���9��T��Ѭb�
��c;f�3*>%^�	���Liw�t9���)���eH�t���D�03<�4#ֽ~�D�JG��iS��P���q��`�6��yEYΨ�/Y�~L\,���[�q��_=�i���-���R�O�D�Z��a$ �� _�ٚ�l��k�ը�ٗi޺%o΀|�N��e���Ƿ����so�o���ӣ#%`���"��c6��X,F	��븼��*��?ZyVrx�����NNNn|��޳�J����w��%����9�l���]N�RP�Y,c����^�FJ��������wI�<~��jQI[�.}ݬ"y��k�B�M��g����r)�ٷ�n��8o��jL��AEzd얛�@��G�T�s[�
��~������&�@��B��zE��HfY����nǫW�X.��y�l6c�^��hQ�F���cS�\G�M�pvvƿ�w?���ǜ���L�=�����{P%���C��I�)B47
5RAG��>��&3��:T��A#V�lh;���6^�z�j�����+�&vTT%�_C/^���v}���c�5j��	�?�,�ą��"��}e{��9���1�Rц���3d����?��l>�mClH�ж5�F��L�k.�/�;�[Q4M3r��|�]
-`�皻�K?�u�z������r9��<y2�?�٢k;88�v W+ EQpxxH�D�躖���1�$�4�ۮ�3G�ٔq(���2�q!Fc��1Ħ���:Z��ڭ�^��a���(��g�F�og �j��5F	�O�e9�U��O�Q����URu]ߨ��3l����T���1��u�͆�,_C ~{���m�
���c��gϞ��9�g/�!�����0�`��`"Q+�S����I�����91��V.z�`%K��%����h�c h���l�k:�`L�EQ7��5�5L:��b68}�MDd�V��7u����U����:ɹ��z$���d��63dY���1��y��[C^��yI���w��c7:|o�K}�����wk��g����T|xn�i����'�s�{�= qT_�z5�iV���@~ѿ�$u�!�%���,�'��!z�vsE�����bD�{�k3�&�6�=m���4eI�ACZo�Z�ױi�X҅���,{�Ӗ�Dxxg����wYU��tƒ��T���״&ݻwoD��-���!b���$�O�~�������n���n�b����HJ���M���iޯ��?�E��g�=�vOhۖ��3�;2�rK���x��W�&IC"���\z1�yyC[��܌�3�#��[�!���,�r��$�#�8g�rK���}�j�BO`z��a7���C~*=-f��,�XT)-�.!�m��5�> ���b�YƤkS�{����ϖ,���������3N_��nT�� Lc�o��eY�/{��%��1�Hc��4h��x��c:��N�8���j��}ey�>�I_�m��)]�m?�R�u�޽���GD1�gC�)5dYJ/�!��������� d����%��:x���	�W�{�5��j).
���������;��[o�r�N�68c��g���*1�[�H�~�P�sb�cg����־#���AlBp}M�ZK�&h}�\���V+b��e9:�������Y}gߜ����AJ��u�j��$��#f�� &B�l�:IKB��Dl/�# mDTq��ӴhD��p�<�)
�ҡ}1I�4|v�&�@�j|��f�Q�@mWՃ����yۊ���;������]�α\���}�sBӱ^�i뚮kGt�,Kf�YB�eH�����Pۓ�]�s���#�=zD�~��r~�v�����g-7Rh���;{�y�o
{LQc%���v���?��?#��f��
�<����ؓyz��ƨ���\B�CHE^�md��b���{�r�d>���l��j��wt�����	t���JK�F|װ�l��ի�^���jeڶ�U�1�"���ߴ�s��|�~�w7\]�����H�zo��ŝqR>>~��<~���7�?~<��?��c�裏n��<~������e�gv��a�QA�(j��w;ޑs.q�4N�p�T4L�餚���Ӷ�f<M�0\�N߳\.������|�ޚ��#Qގ�M�9Mͼs��y�"���b��w-�'�*��Q�ۤYB���GQ�HJ��Mڐy��?y~�PcZ�1��ƪ����rpp���)�|��NO	�ë%F����!t�\��؃[����::����\ڷa�{c��n����,���p��14�=��9UUqpp���!��h������5l�[�O��y���;w���rvv����&��%�J�e@�Ҽq߬S�M۔�2�wH�W�/�N��S�n�������l���Ÿ~ܤ8��=}(�@��8��n�_Z�25cb$�@�<p}?lgm�������W�5��2c9_pz�k3|�QgK���n|������y��v>�}�C�1���U]7��fS���Yu���V�������ݝ�鳏?���9|��G�������g������Ţ��=~�<~�8�'�m���u�e�������Ν;���ivQ��|����޽��������#��n��_�f�7���Ǯ[�_��?��r=�1�g���V�7��3�ϯ���.OO�Ν;������?��G������ӷ[�c�\z��0�p��(��Sq�����S��w���$N�3gpʦQ��Ѿ��n��e��'��T�,#�k=-#Bf�3�Y��2�K���]AL�!����	��Ȋg,wf��CUU l�k6�Mӌ�l6�ZKUU|�;����1��?�)?��QB�/m$�X��M\f!f�eNQdI�y�0i��.������9g�HS
9fdƎ�5�Z��1�W.c��sxx���]�,��
1���eM۶l6..V\^^��/�dl6>������y�=e1c�7c �x}f�Q�o�������`{�k���A�|>�9w#m;Eꦭ�Pձ�p<�1]ō�6#�eΠ}�zP'X����u�n�����ݎYYrtr¼�(r�s�*X.�{�=�+	��{���Xجa�3�����m�H�F��2�vm;8n��X�t�ģ��Є�;u�y��k��(�J��y/��$���h�����;��]8(�͂�My8߬����Y�i��E�m�����D���_�W�a��޺��f;��J8V;�{U����q	pڿn>��O���v'�[���Ƥ)�F����ٳ5����QY�f������w�Т�,�F �ЃI�]��֫PF]Gs$&�F#b�.�5�|�
�nr5}�J�h�0qI�,�vW����m��*)v;�c�U�pJ���C�u����#��>����sk��ιxvv�
�z�O:�R��h4�)�u�:��ؠw�����N^�IL��i�����������,˘�f8�n�o�F��}�q�\������kS�}P��T�������(����w��x��W�%˃��,�ˤ���|NUU��\�s~~�f�D�w�y��}�s��~�{��s>�O���3��Qr��V�^Ƈ4S�%���0:g_E��m68}��5���!��Jz�\Qi[�v[���Rf�jVb���9稪*��B��[�&İ$#xO�D�6�B�Gc���.��!�?�O��ǜ�]�HUUt݊B���f����&��w�E6� E1��5M3�]��ƈ���m[��-����|>MӼ6��E#���=X�4]�y�(�����G���{������#>|HY�����](�G�wPv��H�O�I4��Ū+=�_Ί��6Կ=��e�Uӡ�klB�ľ7�ZQ5ǉL�ƴ�Ĉq�U���(�5;1�V�.��F3+f'��,l4���D$X$8�A��UT�ݖ���HMl���hT5A4�5�v���fp�ҸZb�]yﵫ�0""b�����I�D]�z�g��%���:2o�ع�Bv���D�Js�p�!*�TH�M���K�F��f����fM�	Ar

�QP0N�yI�1I���9�s��U9���LͽJ�.S��Nb���Zڶ�9��J����=[����a������M��VN��ё�"��,DAMT�FUׇ݃ߵG��S?"y�KS$�3?�|��fLqu�'�_��5��?o�*+��kz��?��M��(�N�(o� d?�<=����FUӁo��E�ݝ�7���s~[��mc��ɞ�����3�#|	�-�kgJ(X_]1�9��9!��6\]mȲb��ʲ��|���]NNN��"��("4!�-(燨ɩ�m�qx�./_>��/���w����٫Wx�R��m��&�,�y�j�Z�?}�_1lR	Ŋ�3�!@����ޝy�Swqԥ�+����|�٤Pe�������]ץ���yY�u���"��(�˄��,G�py�e�kX�.���e�Г��o���Ֆ���@3Ќ��gcZm�b����.r$�<U�����%v���u�r?/g���̩��N�����N�������~�/׎H�n�%[��Z��x�#�y����� ��M��#%$�4���f@���������~����srr�Ç9::��@w:{y��t����Z�+�]�|���a��h�]�_^#���
11���FL��J��0b�11m���9uY�5Q�!Hf]$�Iʈ��� ���!�����3E�r�X���8��:&ؠѢ*�˽�]�dY^;��!�1b��ykmK:�`�M�mTTՅ]�cn6������	��jUc����D��ֹ����NUQQ�>�����i%5� jhDE�u��X[���:5]1�N���}�e;��Řh1�d�S���Ҫ��l��Ζ&���Wͮ�;;<�7�9�!�+3��u�e6k�j���������~�O�������5�o�@*Q��bT@}*ݠ@�I���.^ב���i����y�/B���T�'nH�"���Q�e��iï7u���OӖ"B��d8[�1�O#�%x� �A�\ˮlYg;|��
�g��W��@W̉\9Ǹ�g�Ny��W���6qآoA������1Ό±�9�.	['_������&��S�N�I��E$z��M�qxxȼ�06m�����n����kܮN�]V���'-Mo�\*r���W�����9����?����S�#��+���!�v����e�t*{P`��o�1Ӵ�4 ����o��:�y���c�n���!������ܽw��?>����|�ᇦm��ߋ/x��)/^�`�ZѶ-�k	a�:ٔ�*�$���ը��V�\�;s�Q�80*��x�J&J@�1�Vq QP��W�8���b��F���	^�rk�WBhQ��q	Ռ��n2K-֥�c�P�N�O��K���Y��5	~�C׷�T���}x}���m���Ö��*
EC$X�(�^�k0�͊�	A����2'�K���D4�BX7Ω�A�s�Q%FED""Qc4.˼F1�]�fm����La��f��k��<8yZh�c�w��3��umϲ,<���{�����������_��g"��r���rG�d�"�D���5Q}��N�0=�yD��?V}��u��7'ؾ�"���h�n*��6$e�#����۾Y���ĩ���O�����"_�l���X��"6-� �q��vӢq��6-�GK�,�f��>v��nP"B9�Q7���1����?pvz�v�P��w���� ��*(�GJ���ucRAI�:d�^$i����$ۍZZ�a���޽�F�e��f�P�%�K�'b�46k�@���X��Ҷ����s�뚑�:�?;�ɧ��{v|t��W�\^\�Q�?A����_���w����3��uh�o�L���4�3�7E�޴���!�5�J�4���;�-��?�GG�ѹL���cUU�m}V�Q��    IDATo��V+�?�ӧO9==e��"Q)\��D������Ԣ���Q;���+T��!*ɿC1Fz=M��Bc����з����j�9q�I�� ��	>`Ħn;�K뗵L�HU���1�nHE�&����±�w�J��1zBPp���*j�WY � E��@�j��XL�R�V��=�c��>!�"XcG�NH���HL���t����� �Gt����::�l�n��� b�GI7
C�X�GU$�2(�f�2���B���lV!F3�nU�s���ф��E�$�>{�������)����ݭ:r���uf�UjF�"����D��V�.���}K�µ0�t�o���C���������L�!��&���^�����42��T[K���,*P��E �@e��l������A#����@���#n1#���y�:�Ѿ3�Ř��9�S^�x���Wt��g�o8��̐;��\oi6M�v[|r�l����ٵ!�lL����}�o��9�s||�G?�pQQ�9���ټ�	�7+�%	}A�DM�I��ƞ�\Q�I��NB�EQ��S��� �H`����=��v[z�� �n�՛�~���?�toJ����Lm��,"c����>��C�����w��l��IloBTӶ����l����'=�a�z�S�����;���l"�b��R1�1���1!
1$�I�������1d�%�=�!ɤ%~VD�`\r$UQ�e�z�'��R�y�6��x]U%�y��\U�_�3Ϡ��0��u)#��<;�����۶��U�����`��%.'�]ZK��I��7�6�X,��QK�$�.l/�o��q�#���)H�#�Y�3 bDpVȲM�o��\���.#�G�;��NRp��Q�U���,���{Z�Z#�m���A�U��E�a��hu���+˟֮�������ӧ�[:}���j)")�TS�a��`H�nzw���+��_r��|����x����}�E��@D�O�����ЫwHߛ9��ocS����׶m����kG'�<z�}��>�Ō���2�ȋ
QC|�ֲ���5D�����8�XɈ�ӵ����W/h}ǃ{w��J���\UE�#�~_ץ��r��pq~I]��e�s��"�or�n8Q!@�c���~�*����C���!�������O?O)h���;��T9]w[ʲ�����y�3����w?`u���┋�s�֗d�cy0g�I���t��;{g_bӖk��=;Ӟ�S�ox̀N����5d���b>���������k��k�����t�3޷�Xʲd���牎�bS�D�P��mi�Ժ�w͘�v�Z4ڸyTET1�H�;�H�{G��A��W��(�'��[*����c�b��J:N�-�mI-!&D��_�D�5t����~t�Āok����it&�Q��?ט�®k'1F�bUN�<!v�TK�54J�:U�ś���8:"VA=�D�+0N� #DA%�XR����)�� X�I�u$��78k��tmHWbr��]K�Y֑4�u�6uhR�wl-bL:�oO��ɜ��Ǯ�|��I�y!�*bT����w�l�\)aU��s��r+�om�:@��,�����)G=���kT�!�����GNÄ3��k��-������<��S6���/�h�vTr��6]0~�׿������q�&Du���E�&�����8>L���ܻ�٬�{��1�.ru����n���1� ��$+`�`l���F�6Pf����.M�c^��+��^^D�4��l`躖�z�sx<EiF��� ��oZ�n��z����b�����<x���lF]�\\\pyy�u2rc$(h ��������'M��b�ɝ��*��O?��?������uMYe,����e�o䝳�m������q��=�{�f!���k��s��y2���s�ݻ�ݻw��Ί�ԫ�+��ù$�rqq������zX���Eǖ�0r�� �wF�	����9푿069� ����8�O��Ǻ����9@��e�	!v�~�!�{��:���@�u����@Q��5�O�FDL�H�9Bp=Zx���'�SJYBķ���x�1gm��r+1�H��!���&�`�D� ���1��D18��N!`A#���TH� "�9m����}.K��	tɡU�RA��)���c
:�4u��E���֊��k%7^M���/L���Q�u�uB�l[U���?��?2�J��_FUU,���TS����熿���q����.�}��#��Y$��$�v�t{��	��y�o����z��u�:1s���brH��~���y�	�w���T��\�k74�������@���=����X�E�`1�ٻι\����3�N_a�b�z�d�Źl,�0���dGׅ~&�/��u���c����}��Im	����n���+v�K|h0ɲ�5}Sy��Al��+˄V��Md����%WW�\\�%�2"w��a6/��¤#���;�~g�m�Uy�c6��Z��9���,�>}�ڸ��}�ћ~k�(�N���u�f��x�����L4�>C!�o78�]�h!/��~D�i4�E���2K)M��b{dӆ�'�T�Oȓ:))c!��	�A=��	�2V1�@��X0=�-e"ҹB��H܀��y�-�әQ=F!�*�IB �"!^#i`ȝE5��U�I�T$�J������Q^��Ū>C�������t�1H���}��ͮ{���5�K�֌���ǙaL��#y��|O�a_Je��з���H��ش��kE�����Jg��$D/Y���mp�ʖ!/Y�����:��<���5�}OU4�$���]#}İ����_w��& �O�������ސ�"���*��_��6ٴ
z��~]�0��ZF���@��lVr||ܣUk�f�fs�z����ݶy^bm�t�&E�=�Y�!:��i��*�(E&, v����ӗϙ�f=R��;c��'�f.Oܕ��ӵ1��L�;֙����q���+�>U�����������2�I��Jfe����w��O�h��̲Z�X.�TU�ԑe�횧Ϟpyy�'�|�j���'�����(R�|6+�w���:}?�9���X���~��Mg:�c�Z�l6��ݻ<z��}��k��ӷ>Ӡ�,˱��v�5+<x@��R������ *�H�ԗ� U%�^���`�s%#CA��%�D�����ñ�Z))%���(�Ӎ�؀s}#��WC���Dm����������'��W���i�����G�ff�Q ����%R�Qz~�D�I{p������{��m�
Ltt�?ǌ]� �$���\WYw��Y���E<��8��~��)�Z3:s��er�D`�X }�i�����?�8��EY�g�o�.���&��eծ(�:������ό��Y?�����ٟ�ٟ�.���J�ʕ�]�ԵA]Gɦ�r"��Ut1pqq��ppp����3��,�����7#�c����!�?��2�h�%�6�T�c:B�ݘ�S"���5�]�I�_�1=���M%ZTu�쫪��t� :�~��qkR���Q�9�W+�(����%.�8>>�Y5�C�����wPu�OgO�c�h�1Ĥ>ف.M~c0�al�n� �:�EL�䁮k�tI�uc:��̲↰��F��K�Ǜ��B=���BE1Z�S�i�bT8樷��`��eX�"��C���6,fs�Y���9�����k./ϰ�p�H���}�v[lY�-mӄ?<ZR��M����sv�WW���윧/�\�J��|A{��/W4u��Q�a;�qii�qBQt�c(ˊ]�b߀$O�����_{H�"��T�)�2U�)�Iʹ�'�4`5"�������5��N����]���ã9���E�'F!XG;���?��c|�l�5E�H᫳s��/ħ?��������n��a��k2�:�.8t;d�
�{�*�n:Z�Ĭ�n���G�*@�$D�د�W��:O3o�m���_.���Ͽ]�T�U��w��?����:Y;��h8;����o�#%��-&z�A�T2:brB�W[	X"&v=��}�,K���m��|��/^��,��ΑYG�8C�
�،�_����U��bA����1<z��|N�u���s������%���ylϰk����(�T�d�X���Z���+}���T��y�5[�U��!
��d����wԈo"�$U��H�q"i�	�����z7�A�92w���t��9�~����+f�*Q2d�&��@�Ћ��y��ډ)Ö�*� �'t�=��������_ЈnS�u�	�"�Nh��8�n�g�q��0M��7,Ĩ��WW����t7)*!]{Rv�ZK�K��&b5�������|kC��4�3b�X�����U�y��*ۧ�=��;���=�����r+���͑9�sng�e��7�?4ָ���bq������ܫr||�n��'?�	>('''��?��Ç|�;�[��ЦJ����f��>8'�A%r-r�����O�"���(�V+f����5a̶mS˜/5C��uUUq|rw��l��5�1de��b4�yvcQ��&UI6)�����4"�FޚI�J}z��K	��!��}&�]��6p=��sT���O�<��'ed�&n��Ʊ�D�e4�TM�׹a���cK2#��>����3^�xE�4x�l�B��������w�4���PM��Wu�SN����N��i����yV�>��qyy�RB:�$F�r>C$����~AA7�o;DW��PsN�v�<u�i�@��fGizD3"�6�a~��:���s���v|g�1%����D*�jO��:ƧGTԠ�;���Ħ=�m�)��(s��Q�A�y�ٰ�6��f��?E����}$i���ck�A��իWq��=���z̦
�r,�����M��6���qy�bWo��u�����9�>*1�^��5�RV�Y�o�njb���Y�(1�� kՈ�h�k��"j�ب�ֈ�tm�����.�� &b�11F%��Qɫ�'�1VĊ��%&�;l/�"Q�=�$�b�%&R,�ԀŰk�t�%�kɭ%K���m�c��#�!�M�PDERn]DDQcDȋ�!�:��V�h�ѐ�� ����$I���DMH�pbF���(z�F|[L����<ύB�#UQ�n6��ƽ:�l�3���Xt��^��f�uu�Ύ�Pxa�絬Vw�����>4��#w�]��Z,we�>]mοqy1__m���#r�.�͖O>���G~�_�:��[��~�������w����z�n�A�������c�!����u�{|ұy휦��s�7����c888������a���8�
�?R�;�IE>F�(�E���`$�/gE_u1.E$�7�dLS�)e.JP����װ6�C.+�6�kS
q$`kPZ���_��NSb7y	�>��zр�I2���'O>���Ã%��"��K<���#���c�ݎ���� J�yֻ���J"�����iȳ�!Jd�l�ϒ�rQlv�XU�/*��6�!�(��Sn�v���oB��3�����QV�jFQ$��#��A�+m͚t]c��a��u��imC�4dE��{��]��A^���Y{6��*q�G*�TO]�~�_�x�u��&�� �o�}�:1�����}u���LE{�A�����{1��!D%(X�1�r�9�����;	���ϟ��:!���z�}��^r#��0�^��NM�ӛ��m[��i��w�����GwX,c����fKV�D�]s�WWk�THB��qآ����A��^�Q5Zkk���ͮ �!Q�Zc%`�F#.�P�J�(i�S�F�� �ص�c0BT�h�E�ɜD��x�,��Q5	8%WL�Iu&����h��|L� �C�EoQE���C�ƣbS����'jp��bTo���Mu&����D5Q�(*&`Ԩ���^�DT����A%�:qV%D4L�����de~EP�ZŪQk�$�K^[P0Q��D�"����Z�}�pyV�l�n�?���ؼ��mk/W]4��ZSΗ/c>mB7��;5���ms�`S>}��r�f��ɬ)K[:g�u}L��ϖ������<���'���<����������~���<�麎��'�>�����z���:���uz��N�x����nJo��m�ޘ��}����X,������v��7:H{�Q�+�-�_�xfՒ�,8>>����fC�J拜��M��(g乣���,+0&�cL�Ve(�W�}$���e��-ƪ����[���q�y�˗�	[;�\��'H��p�wbBHZR���4u��O��η��-֤��(�4�6�����Ǯ�����$�@S�l�[ !�yVpxxؿޓg���<{���nGY���'�P䡿�~AE�1-L�˷�o߯!�r��}�/ƈW?��%)�Sf�;ܻw��|�^I{y�Q��a�|��{]��g4�ѣ1`p�����C�1�Vk�.׈���)���>�W��x���_�o�&"��篻��M��N���J����zA���j̐�����$g/�ɆÚ��ڶc)ˊ�G����|�;����=�����m9??�B��m^s��Nݾ�K����hc��Q�%�Yjƺ^�YoJ\Vp��{#��g�~���Ϲ�����紭��k|�gs�>�2#sE��U��,�X۱\΂�U\�bи���^Y�M����T7�1DDB�k'-5�0FZ�N{�R�bD��a��B�@�E�5�5�1#�%CU����Pi���AU� q�gD�H�C0�#ј$ *�l>����(��b�H!ΡN�LP�1�^@}J��֤�a4J��	"*B��Q�`� N�1"bzb���+`D,j��DL�1F��g8��N,N}aqI�P%KM݂�(Ɗ:�PE��'bTd���fWKS7��U��Qe���(��b��˳�6��6N�%&����]G��p���s�x������ӟ}2����Kg������~���{�71��gO������}�v�e�M�^�I����h�D�b5L~��Z�q��d������ hŵlF{�s粛|���A����������ײ�J����s��E��Lf��UE�%�n $j`�p0���x$�dO�T4�&6jJ���p�$��b���.����ͽ�t��`�}�7^4� �ɬ\���⶧�ͷ��ַn0M��@)�T->b��������.ZB�hm�T��+}�) A��(���ֈ�dD1ZU
4Zg,�e,��-m;�,�<xt��>��O�;Z�9��mFw~�2�G�a�m��Dƌ�(�x\���Ÿu�![Qr�y�eͣ����{�wSd1J�6��~���8����+{W�&��O�N��2V꬧!(|!����>x:��u��ǆ�A�0�%� xK�v�g̦�NC0jz!P"�$G*�	��{0���+��'�8<�zL�^ 2�E��2�H���4�?�'�'p�B�X,z��k�������Z��{~�q/<���v@��٘[�������+/�ҍk�l�@5�'�Gg.���m�6ı�8E"=?�u%��r���w�]i��<�gP�Q|����G�q����Ѡ�!u��>����k����1� ��D+��4@�_�&�"w&�m[;em3v��V���^�_B�6�(�\���>�Wo��V�g���Yk��+Wx�߿_ ܾ}[������Z��U�:(YԕX�ЎGE8���s�oo/���$(��tz �U5Q(
?j�6.di��ɲ�g��"`!4!�U"���ZP�NL�MJ��B�.Z' M�S*(+$�SBy��RBz/�tN� B�
1�/�`��2�XQ���B�P�F���gI0��R���)8�C0ʃBH!\�W�hB�Z��,=ai�.�M����BdƁ�o}pn[y�-�HJ���/��?F΅�y��;����_�B(u�>n��_�u��ڰ�f����2�����)^=?<���ի�x���������ʫׯ�����{�QU����5��M��Y,�H\�|�B�8�Z5U���J�I&� ��K���F�ןdu�P;-)D�o����J�_�.��9�~�u^}� �و�i��ڢ�sF����Ƶ����m��^"�    IDAT� *�B$8�d�s1��\ܬk��1�B�ՆJ�h]P/�@�#���ݽFg����c)�M�W��HV7"�
8p�&GQd���5��ªRQ5��%�t����X�4zW�Z+�Zi,	�zpF)�(��Ҷ�Q&��<�E{~&�1L�'N��1O�6@w���Ma���ה�EN%B�vL!X�*^�Qn��,�~�C}��(F�gG�h�����
�c��,/O'�����i�,�9���g)W��{��	����OJy������Y���_�����$?X�V�����X����]<FE�	R��d��ǝW�ɛ��;ܼv����іs�Y�q�ڵ�/n��|�����K�,˲��:ڄ��f\�������S/k���9|t�|�$7��tʍ�n�IE��`c�U��ٔ�h«�ޡm]�&����> Bt�t1>��/*����k�e+�:w���xY��g�TgR7�1b�_+���?�hƍ�r����]k�r~|,D��HQ��9���^-��΋�B�\V2m��cW�4���u�T"����)��-N1*8畲2H��W6x)�t��ޏ��FFI�*��J
�#��ҝ�,BK��I�U7¤V��A��R���U\�Q¨�DV�m��C��؂���5%����F{-D� ����+�Xu�C���<���uP�U��B@�&_��̜��if'�X��ű��+j�r��F�Vu�װƸ�mE���kN�3�PB0��6-c����@cãr��>��A�X,�G#����{�'2����2�̨�^��7�1�����?�?�z��M������X�i������,�������'Ҷm ̲��֯G9��'��l�N�?�#ȡد�'R1*��)�.�g�c4s����]��|>g<�!��F�1�;�ؖ���oq��mv�v{Ep�c�"���f��%8h��
�k-���UJe��q!2B"���{WnrkQ������}C��U���K��1[�X����ȁ�9�q�t�WcGJ	JS�%mk�.���A�<� (�̠���-��($BE��YI��
���Oi�$��e�/�VI�j��l^�x\��ƛ�� b͐�Q;�6���5�[�R��_i%vV�(YAH�X���ɶ!+[[[�y��������5��3�v<YW f�f�R�8E!E�۶e>��|ޯ-Ҝ�m��o�6�Vr�خSB��I���u�D��	�0���d��yԾl,m3����5����������F�&h�|���	����h�����b:����#|�}���)�{�"�3E1��O�� �m9:=c2��d@*���q1fk:cgo��x���uՀִHB�≕�A(���U�B��Y��A��Ω��_����:�3�te�e5,��$xӜ��4AklfDH)d�/��Zj���Ef����J���@��"ӍkE�&���a<��E��)R/3��v��j��Y�V���@.sh��Ω��ZZ�h\���-弆�	x��m0~�۶�ң��^kC�
�@�(*x�ڊ�P�IW*�t-���!����I�*���RZ��.SN���{�H���VZ�s�\ȫ��:hmCM.�R�;���0˰�b������ ȂZ[8�E봒N�����a��c�\:)�h�H��U���L_׳Ҷ���I���K��;�^{|�Xܽ{��J��G?�Q>�N3�n�\���rY���ٱ?��l�_�1j*W��_��)u����X.z~C�XQ�2M�E;;;��k^~�����<��h��4��HD��r	��y=O^��}�(Ek��ҥQ�aX#�h�h4ekk�K	[��QV�%�Ķ2EV d�m%M6�s,DId~;�]k,��Ź��ֱ-�{6u���"���qaPz���
�٬O5A_�f��ջ�HY��6�d:�!�+c:�,��ei0&��Ľ���n)�U��K��B�|�]4Yu��-&K�K�Sb	���*�?3�S��9pP�L�	����Ǉs#�>���n��,��0�8�r���n�x����Ŀ�d�w�L�� e���-n߾�1�b�c�X�����x�J� �{�(@/d)힎x���_Ş���W���"�08M�(놲�T����P�e���y�[,��|�f��b�7��f$=�yyv���H)���fgg�=�1>�ivv�z��ml��-�A�0�c<˘Lf��cw���-������z�eEU5̗͠i���ŕ���|o�ʃb�5���ն�vP�� ��(U���i�?��?�������cl�?��?6;wv�ݻ��ܽ{W�+�<�n������ �O���uM.��\	������t��6���ݻ]�6'�����׹�=���x�Aw�#���Wu��c����R�E&��t\�Z��w�����?.r9j��s����3ᔒ8ȥ�Rz�XN�B��.ŸiJi�N6۪�B�|ڢʕ��m_��p�p2/r�Î��K9�b\
�j4
EY�J� ��U= ��)�쁗R�u�hfM>�TB7e��,ggJim�k������'����ޘ�F����\iSN5��,F�O����������m;���G//���GcJ�+H�ܽ{W�����d0�a���r^~����'ׯ�����>0����-�,ʒ�|�U���M�s�jٮyI)
�@댋�9R(��":aܺ�{04䞥��1�:���0z5|]zm���E%���W1���Sc)�u��L%�Uu��/*&�	{{{��N�\�}/Ҷ-{y��,;���`�i���S��PJvi�mO;;�loo��k�`kg�E9G����ׯ_痿��ZK����o������X���mۧL��y��F�NJ�X�1������$:�$���R��D>����,K�g�ϳL�#B�8_��5e:����`��6F�mF��W=؊Q�؆-I!%�d=�������4ϴ����*Z����I��4Q�l8��s��z�F1.2Dp|���<|������_�¨JȾ��t�s�\L��0�IU-���f:�0�a>?gR�}1E����%���B�P&R���ӚϺ~�⡽��l����阓cz�t�P�uEX�������G9]������ �4���.:��PUι^�nx^J���";U��c�ұ��k0�B)�K����4���E�W%R����svr�������7پ��:fY�F�ؼ��>����`r4�a�����O�1,�U_����˪{�h\�ل��bL�:>��I�����ߋ� BD�����j:۲U]����Z�N-����]�����O�n�S�4h{�O��O�B�w���@�v/ ��Y�ON3�d��u����������~��B�&=��m��+���������w�>����+ ~�_��O�I,����],�)�O~�Ez�}��������L:�&*��O��Z�{>�������&��𘦶\,TU��m�;⻖Q�$6�o��|�����kO�mگ�n����Sۜ��	C��&l�� V��H�nBNN����ϱ6�����9:�(��l���6�ٌ�h��2�R,�K�m�P�5��ؑAJ�Σ��ry�w-R�.*�N"�lo]�ڵk(ex3�,�"���׫v������o$��1%�V��R��r�����Bj�#:N��zK]5ض霅�P;nd�g�e<)�(���K׹ru�,����d���y�8���
NRt,�x��k��;<ݵ�a��%i�]8R����cGGG�����7��|��(-E?߅ E�dq.���>(|�B���_�E>��
]�Pֹ��]�>ϲ�R����v��5�N��Y����&��4PI�V���Ǯ
�E�s��+_�KW@V)��CXkeY�<���ixmdX�nױ��#�Jc1���,��w6��9#��"���T�1|>}��a�.!��j���%:�v����\\,8?��kAz]��Z�������y�|hl0:ڹ ���8/���_�n�W�~@�W�$!�B����֜R���-F���%�V���1.+���B5ֲ\V]��AL�@�GLR4 .�q�{��;�Х�:5!e�_�S ��FA��{��D�u2�����_l��%1�+�)���,�Ƈ�׋q���R6Q|��M��Fi��He]!����a���=�HK�u�tE�E�G)cd*h���J��/�~��n���x�=ί���s�]��@��$>�F	���qH�2����<x�����s� :��ὥi,�q�2B!�Qp��0N��0��(2ʺ�:��b�G/,� ��qL�&�(��]�$��b�/����>��s`�s!m:m�2?�`~~A]V�F�ј�Hk�u՝k�c�Z�4-��<Q�5˺BJ:0+x�]����Ż�������_w��߄םM������5m��@��C��/�����#|��E)Z���!��Tb6F�2��z:~���] 9 p��o�RA�R��i�
! ���T��s4�C�6ri۶����~s�F��OT����'���:3��BPwm���$�_�٬�gi[��%U�62��U:����J��"�`�Rʠ��� ��r#+����}/g/�͸�A�*쎔z�;ޮ.�j�[��L+#�m+�Hmc����������lş��DN�[�l����I�䋤��퐿�*��b��~���փ�T��-;u]����5��x��A�Q�͒�ىo��ki����L_���x!�"D�hO��-	�&��E����c��l_٢�� VU�_�H<�L���bY ��u�x}%��9QH�-����Z"�Ƈ��A'�#�z�T���-R	��<2�6EⳮsN���{R��E->(�Δn��v��0ґ����&�֚<���۷oRU�pzzJ�ƴ���IN�2nܸ�h4�������DG��� ���N�`�S�C:F����Ն@-X�C���k���4��}l}:�����f�Kkݧ8S����UJQ5yV :�<:F���YA��H�P]z�B�tp��^?��2��>��-���N�B�H-�
�����n.|X�9���t,�
�aT3=��J�h��&�7=��)%]���|�|�<�i�lL\o�~J�a#0M=uE,8�b����� �B�B �]�7��_�	��F�Aߏ~����VB���k�Dx�\��M��=��r_�QMc�VBi���	��������,k�]!GU�4sXq�I�O���G�@�u���@_��z�=/�K��fD#mr)�eQ~"�z�`a�֚z (�x۠��f~qF]��#9wTh�rk�t���"dL��`l�-K�����N��Y����ՂE9�n+���X-�k8���_F�R�\�0W�ù(vj�AI�:���}l�����،<�jg��w9*ʾ��Z�����=v�jI���`��ԇX�m��M;���"I�Em �}#���j���#¡K��o ������tʝ[���%�lo��3�Q#D�f��7n�e�>���������n��R�i^��|���xM�9̗��Cp�����ۜ�B�\nC��#
<��k�ް7y_������ZO�bb�4�d�QD�*��*���يk����f�A/���E��#GXE�D !Bt���*��!F�Et&����ԋ<��t�����Ɇ�z��4�ctUB,KiݢXU�6�W�~Ew��ή�����>:G���7"/�pa�r��Ʌ_�WԞ����?V��Z�L�Z_�PI�}�loX/F���!h��Bʖ�jp6V<�e�b�`�\R՝j�`���gll��GEV�6A��ؐ��;������nO�����i#}����HBFmom��=��~d�8P�Kc����bR�T� c�B�ض�#��n,ZOb@Į�6�M`Q-�M��W�%ی��Q���۟됬�eYWuk�wR+��նu(�P�'ޢ�D�碦_��v�z�.��c�g�/5tH6������ �����(� 6\�s���d?�g����lm��ٙ"$�&S�� XJ�u[��LF�Q��� o-Ai:l�G�DQ��:ܠsI�δQ��˾�%�>R�v��xX���@k�^d��=+z��J`��[�	!8??,0��%�p;	��<��{�W^����N�^k&�(g"%k�����A���`�\������w���i�}���k���/t�͡�v��m*lS�J��º��u�2'{�;j��s3���M��a�_j����>��|�9�v�AV?��c��N1B���]1�s�{'D����E&�pA��?Uw��w����ϔ���i���K/�d\��ڦ�i�ۡ�oi����1�MdB(B`�����CU�,�Kʲ�i�ޫ��L<y<��|��RR$.ti�4!C���K��~ÈFz���5ӂ7��t7��K3D�	�u�5Z!B����M�S��6ѳ�]�^A���m� d�<�9��6t���bU�`p�%�g(=[Z���]����^>�^k����09L������%�R ��?�w��9�[���g��l�z���k+����Jhvw�0�ls~�����z�!���b��m�@a�jx�C`ӟS�u�����'�c�|So�����
@�llϩ���{7�1���w��Z�CL��h����G�M���	e��;��u�����Zں�>?g2ʘ��\\��qqq�����8��iKU̻��ܹs��7o2�N{�����J�����G�qxx�GĆ��i6��Y�q��-^�u���h۶�qxx�9L�OgyT�t!T�'&�-��*�����ʕ+loψ}������dru�9��!��߿߯ǩ:XJ�Gע|�YbZ4�@�,MS�45F\���՘N���4�W�<U�.պN�H�~e�������}�C)���	K��&�)rYe�g7�v��<���  ����',�K)�T!��)������e���!{&����Ea��B�.��M����ŭ��!d.�Y�ڶM�P5�Wl�4\\\pvv�"��{z<���a�b�e�͎+/h)�>L�$]�M�aU`\��?p��TBpx�ҴqS2]�!.Tݿ������RH���xD�F����Wd��Z���ֶ����9εa�F��Ǐ���REj:ס7/���d����{\��G9��]�"���=����X�� ���Ǳ�(&�|�\�r�G���s||�Ėa�'�6��#+_�ml�������z����*��}��� EH2u�I��X�y��}�1����y5M#[ư\�,�
�$����(u^r�:����=><�(88�k�"�D���d���-i����|�����7�d{{���^$�/�ܿ�w�}�>����}���Z���lM�N������?����e���>�������=g3����&r�V�h�x<�ڵkloﲻ{��l�U[�uG*��6!B�Fݤ��L�yN�\a�!�/Yn4-�֦}�Ź����=�6#�J���x=7��%o���=���E�}��5]���22����{��%�u��g�Dk[��D�TȂ�)�wNxB�k�����X��'?�r{H_ۯ͞�*���ۚ��Bη��(������C�~{g�:[�mB�z�y�E����t���#����JM��Y�e����u֥Z��fк���NF�U�}3B2�`]����)�#P*0�Bȼ����2��N@+R{-O� H�!r�\@���Œ�j�"�;�"�׫���=��#�ж+1X����N��B#��X�AZpb��;hs��\ń	�Y�-1£q=A^"A��;!��b��"����Ł�ӿ��T�W@ ױSIE�5����,>�m^�l^st���6�RKPc��tdN2��A��l���.g瞳������;�!M�rxx�T�(�4
)A����Z�l�2�Rh$���8�dΣZK)v���b
�G��GT�#\3c>o�׊2LX�#=N7�� L�h�/tu���ʣĂ�{���������	/����#>�茪�bUMۖ]1��i���S�F���A�!	,|p�#>��N��ͮI�1ʵ0Q�i�αl�����Z�Lf����    IDAT�r=XQ�l�����a[a/.x��}�|��5|��G=�mK\��"$�o�^�oα����(�>�����!o����(]����t�W9e�
��h��#�2
�y�o3����_��w�-����_B�d�s�&к@���AP7'y6��+���0�����{�G���y��QL����¤�c����O��ã{d��)Y��i�[��	�;Zo1�m|0\�im9)+�|IiA�]\�chj�4[ܣ�-�y�#���-M�E�����O??���9���x K���K�+32���~YU���HtW���Q���Zl� dF��ف�ʠZZ	��u�[]�%��p_J�Q�d2YE���W��L�3�`�$؊Q����Z���m��]�gu�PE+����'~���5��v���O~�g���F���e�������m4��mS�m���qV�\ۚ�r1�"!hk�H�ZY������t��S}2��i���<~��'m:�M��I\�gِ?L$sί���+%k �@7��--"��I��e�����ަ���8Kq\���pzz���9��"�r�_�o�w�R�[[[L&ڶ���,VC�RA�-u]�eLM��]pzz
�����t� �F�u9�1)
����0jZ���c�2X�%��R�bDEM[u�4��9??���ggg�(t@
�)�e>,UU�ӟ����^��������^A$���\�� �Eɣ�c�j%>�9�6��Y��_�6]���1J����*I)�N�YN]�#���>���G9���|�"�D�n[�f������(i�9�~x�G�c�Y$��UJ!t�����9;;�W_����=�����ƭ[�\����"�
�����ߡiJ��k���=���lW*�aEt����޵\�ٍ�����&�=�;WؙL�'/���n8<<���}���p���b�������et��O�~}�1��dC�4����&��2��g�&�h���v~}�4������<?�=��lD�N!��cc@�	)����Tq�w�{�m[?Q�|��ھR�D��o��y�P���������>����y�|欕)%�8��2��I�uC�Y�n��?ib=m�]69�mN���0��<�g|��6�7\��0!�m�I�V����1i��X�f�{��sH��z�*����P'��x�ˈ$!�?����}�������I�t�fdQ�,�cggg�����>GG'�Ŝb�Q6U�Df��޺��JF��8M�s0�C+�4�}C�<��P�������9:9������R��ô/ҵ�ƴ�!����Q/K�}��-B���� ��K�p�tk2��o}�;�nvU����s��d{{�k׮E���'g�<x���t!�����4K �����~CmMc�n�m�_ҡ,�`6�f<���t8�y�`������cL�۶�J1.F\ݺ��{�Ř��өb�&�)gg�|Y#��
.��he@)������|�{�����s��U�Q1c
�� I11�~U#��(m����()P�T� ��,�|��'����f3�2(�3ݽwx�o�Z��Ԓ�(�m�g�~�/~��}�q}.ж5�iim���E	I��]˦S�i��� ��5�`����mF�6�线4X9KB���)�����Cǉ}���?�������f1x!;�2!@�y��|�h۶m�.���eO���y�PJ��u���������U�^�u%�i���n�z���3�c�/��I���?)�&�����z�M�˵�ަ'�����=�t�B�����$�O�(wQu'j��V��<�#}�i�=�}�-��C���^�@���0��w����"�z�m�`%��$�?����i��T�����:23��.��f�j���"��j�Nx���6�4��9�E.��0�B�0�I-τ�Zj�.]�,U=_E<dlٖ��>D����j��E9?���u���3<x�Ғ�r���)�����C�b��7�z�:��'a�)�Z+��7\��4�֪`���,�x��Ke�{�TdZ�n������W��/x��88���&G�8}kɌbR����~HӾʕ+c�f��x�W��u��ѽO8�#@�LNn��X/OGl�v���m^z�6W�^�+�r���m\g�D
M�%���w�޴-6x~��_�����xo�ʐ	�ف�����T�9!������l^���j�NNN��_�����?e����;/R,�����p�F�n�t��)�r�7#zC����a�m���y���ק��/�qY�am����sx���ވ.
!�A�����|�*���w��]N�|m_�.}?��G�,)G�r��<7�}k�"ǅ<X[�U�ؾ��m���n5���+B?	����`6'³#}���gġm
i�k�T���&hn�����3-v�h�"�i��7�҂��qn7���'�����)�KH�ٞL���6̛�
��TfB�{���I�%�E��/��<�p��������)Zo���KKY��pq���I<�'�g�<Rx$�Jx�z�s-UY"���Ѻ�T���G����nh��E=%#J�����cQ�?:��.b��!k���2s�_֑̿����������Q*� ]��1�!p��M�wv����{N��D]6�i�g��xo���Z�@��-e���K-�����Dmȶn�R�<��9?��ˇ�>�v���@l��#׆"74����|�U��aRL1f��Uv��"��X+^�4��A*�����[������Ɉl�̜����G�89����n��׸ze�"����o��Q���S>�A�Hap>�Enȵ��Nb�*99:`<���������-���}�O�	�Qt�5�9��E=���#x�Qp�Y%����˂CG/9C'p3�;�5x�|��eA�V�Li�Rq�w\�ZO�򑻙���� �y�k2!��!��}�i/..��/���E��I�>U���fu!��.>��=��R8�2k]�"y�A�tΒw�Ti,�G�6A�����'�U/� ���'�Uz���n�06m<��u6\L�����M��t��ӳi�s��9���@��@����0��#i�)J�e#cG�t�����soC�{��(��>V޸q�o������IPU�Vv������#���� �7�.(��3��F
��l@k�eTu��);�>�(f��k�LJ2[
��)�@����)���T��ց�vR���˷��-B���lmm1G�7�N�������D�.wP�|2f�6l��MkЗݒ�L]V�4�b�����hIP� =���P�������2����Lg�Qڠ�F�����G\�q�7��m�����;c���9����+�������!3���)o~�[ 3�v�dň�_�;�1ϸ��<��n�Jl"���r*DY�kj+�]KSW�u	�#e�ZVZ�L�ZK�mc�8HB����ȠR���:��63J	lmfAV�T�&ْ��Pӵi�����w��a���;��瓢|�<BH����(*� ���]q` ��T��/���9B_�W�}o��vѶ���#��*����Rd��s�;'���d˪�5��R Ն��:�2�7�'EF�'z��ϻ�Ƕy<���_Ԟ�"H^�Uc��_������{~<GÁ7�?6��.Z����>k[��b�m�l'�b[��}J$�U7����k�x2����h���Oxh[�/N��BjW��˯F}�N,7����CzK[/pv̸�L'�MC�ZH�-}A��(+ٽ}qԧd�

.~^��l_A/�,D'D��\�޴iꔢ+�G��ҭ[\�~�����6lmm��=������C>��s>��3���d��R�9PisY�����:g�!1�&�b�O?/|_к�-�Z��#��<S4�pX�"���.�������}˻��:Y�ڠ��z�:CX����;�����?�6W�_�0����'���|��y����G|��4U���n��c<�p���L�S��#ڟ����#��drL$�E���6Ff�%3D'��%���K�H|yD�*�S�&�s�ZE����/��G�9��^�o0��Q�˲O_��n�����@��>����JC:A��د7�!RI%ʵNz��!���l�/tB_�W�}Y�����N��`~h��V��Xj�#B|P���\\�b������ڶ�ҽr����j��\О����_�'�Ӣ|O����MI�.W `��6mC�Q1�.=��=�mr�.��<��y�n�U%o�e���]B`�D��޵έ]��jrP�g�EH0&c:����KU׼���\0�M�_q��+\�v���=��������R�������'L��'��e�s��N�?BG1��zįA�nu\2F���ƬG�AU!�`�V��D�SO��0�DG��U�����:�m�N�r||�2v����ˊ�j(�&�d�b>_P�j��������zd��q����i�T��� |C���%A*>�
���e	�cr���	�~~���9�o]#�69٨��k�|L�O�fʝW��|����=����:��䀏?|�w��w��3*&h3bY9��'ܫlӐ��ֈQ1�(
2}��ͽ�?���1AI��8��5��:���#eҿ��a��a{�T��[,bˌ�}�m)�k׶4my���;�w��	\]f鵛���Vlϲ��!)36�	�9�.=�'�כ�/t��Y�"���
�۶�vޣ��(��J[�6~���EQ!�L��[���·+�h!����9+ j=���Ӯ����p�X�QC	V��4d����~�EC`�xp J�~�%��m��S
�o�tC�LmZz,�K�RvZ������g%��������A|�^j�7Y#D�3��z~IU-㢗�]�2��\�w��	��A�:��$���J�`mۢ�^S�-��@�����W=#��燭�ڶ[ػ��m�RQ��...PJQ��r�7t�x.�%�~�m	��V��ӽI"�1��y�.p�����Y���"j��lw�t�ŽO>�O>A�N�΅���P=??G�t:f�5鮅Z��q�	��xa"N��x��8,�HU�����Ti�e87攎�R3M��ܼy�s��atN���%�~�9�Ucx��7�&����,%�ɬ�F�e�d4��D�X��|K�$�eS�yF��(�춉�i��j�B0Oh��O�E�G�G�@�#�K���$�P�5����!(�b��3&�)��S׎�7n�ƛ�ag�!X�Q�x�d��?x��G��#S#�o�1�L�8?��'q��o�v�I�G 0o*�]��믿�{}���D�ڶ��]d`-!8��h�=�}w���"G"��e�
i����MS�ܬҠ1z[\>+/i���Ul��/��D�e����f�Wi]��Eֆ�9Yz<��9}�����&�iHQH�6�M)�Z��dY���jq���G!��#2���Z�P���t~t�:�����dk�oZ�Fk-�.r���͵{�ry� ʇ@�C|6+�`5���L�o剈u�1�w����O�e��
�o�f�ox�c�*웑���!��;'�I�����t���]��\��7a�]�a�Lj����5Z�l=��&�����w5nW�b� �Ĳc����)3��lo���͛�<ċ�h�sx���~�s�O�;����3�A�B�9 ���)걊\���}!���9o�c�2�qcy���|�7n��g��͛�w���	�n޼ɭ[/���e�zf��8L�{�c�E�%s��n1Ҵrpc$�XI- \��'b�G�G��cB
�A�h�L��B�T��#
d"V�m�x��u�'̗%J��b���t̍�7�y���%! e�ֵ?!�'bJ�!E�:e�+� +P4�Ц5<i�^���q6�6���(CN�e���|2��S��c��K��9��|:.�c$4�5�S}p��,)�����5���F�CX�Z�f&��[o�~�<������������n<��&�����Jd�û�!a�����ZOUU}��չ��5�N�%���$�#V�ڢ�eY/߰\./%s@�	�6%W��>zR�q�zuB���wi߫W���&ppp�sm����s�{�1�F�~[�oӫ^'���6E)ʴj����m܊���;�N��൑��X�9Ej�dy���yUrpp@Ӷ��#~�o�u,l0
k�Rj�2��������+��L&���7�:����<v�H}WS�7i"<{ %෪��w�v/�T�l�M���C...��f\�~���6U���_���l6coo����_�����-�n_����'8��m���XW�����.8l��@J���:"j�I�q��k �Z#�J�,� �֝p�H�Q2�輏�`	�fgg��~�����1_�� i��m$�h��h�k׮��K�����-��(�8օҤH1D �틄�,�c  �߀��W�MD���k_�Ս��_��۳��X~���\]�gR6�POs�7���a��y�e��!(�cr
c���Z��8F��b�M�I!*˼Tm^
{��6��N�Aߵk�dQUҵm!
�mx	P�����&?�%W���ٝ�{>FD�SD&3IV�J]��%Ah@���� �hh)�J�6h!h���$�����Ph4��"����$YIfdL>��fv��{���##��,�ٴ����xG��|�;�q V�ng!�Ty:���V�N�q��"lӃW7f��.rڽ��`a�:)���ӿE�J�Q��?W�����
�?L*C��:\-����͛7{q�rqqA]����_���~���?�n�d|�M�}
���c�o=S7�j���-���s
�v'�!��u�,�8::��F���E�ц���s�3���py��~�9M�k�&�US�i������_��_SE^Q�K��of,����k ���/q*~0��������y��	�����w�]�x�.W��]Ĺ���d�ܦ4UU�u}��1-�َ����c��U��� @�F�"%�^���_�d>M�l��1Ɓz���FR@5����X�'-x�iRpt|���w��Z�� � %vr�|FQ8#����Vc7�`�Ez��S���i=�Ȁ�+=�A�b�%����1FT�L�!����^sJ@<��!�X�D�jp>���N?g��+�p�Z6|��w?wwN���S�]��]���e�����bY�V�1"��k!�x�
���8F���Gu���_��?*l��������hT��2�!�6u��M3�<��@�Ո=���y㺛lhV=M+�P�e�NlW��:-�ˀ��Ŵ@�Ĥ��tLA�"��f���i�X��B_��w۟籧��1�ئ�v [y��Z���)��P�+�v��x!�~�>7};�=���+l���4-��~��|�;X���ϸl\f(\IY��tng�o��&�~�9��4MC���0����t����4�����U����.1�7`��϶��}�����l�S9�T���Y��uC���s~�ӟ1+g�G��b�prr£G���@2f��WdW�]�}zs*ȏ=K6ݗ�N��-�q��&*��v+���5�w�}�b�%���fB*�Qk32���ɞ�e��4g��rA] $�؂���Ѕҹ��_�X�f�%�!�%�;��3 *1.Ukƹ�uC��|����8�y/��@��n ��j���_���]��)�����Q`���l6)/�q[@�2�AMU��i,��u�@|�_{#?~'���=�������;+�2^\�1bct!҃�8.�S[��؀i��*����ލ�v���D�RNۮ C��f��`L?{��/�������_��]a� (�����o�Y,���^�S5d�
��θ.��c��
���������<Ϲ�����t|�(�Y��X@x'��ٕ>�4���3��!}2�]�e��ߧ���}��o����_���ڶe�ڑqN�m
��4?��OY,<=9�k#m�	!�����;�|�q�M���/*�~`ڧL���~:ޏ��r��g    IDAT���x��	�}����T����_>�����9�����o�W�B�qxlH��뒗�`uc�h���'
�k\@�C	
��z���s�L2ж>z�lBǦ��1DI�W1�z�e0)�,��jr6lښB3�v�A�jE���_Ij?*x]NZ���a;g��w�Ok?����1����Ϝ��o��F4��]�igN��]V�y�^���]���_zc�G"PU{�<������Vk��?��˲*���
	�*�JQ	Ƙ׸n��������,�[�.����m+H$�Du�*���T�0�`�Y@w�5��l\���2r�:�D�����rd�՝�q��M�_|���a�ڶM��5�H���m0Nd�
Y�.h�0j_�~�/�x���]�ї���������_'��y���i��, �l^H�W^6~�v�@������[�U��{�ɓ'H/#���O��|����٬��2���&����#BE��%������O?;�Ó�G���/.iZ߳'��נI�f�+�(ڂ����\0�&'��j���10��|�Ij���P�%1��"'ONyzr�r���|NPX�j��dY*�I��  s��$ ����!JL���d�w�o�AVfUNV䈳h��+}��՟!���OQ��,[�B�e�QSg��1�N���^9?_�\%V��cFr��i��3�.3�J��,Q�.D2 uߵ��M@�v-�}fZ@,�f�,I�����B ���#2^������Cfh7�m?�i��1ﶰ���u߱�ױ�S"c�=�}q�����o�믿����׿�m�"BQ��Z�AИGW��ߏ�j��裏����Z��bv�W�q���B����a��M|�Dc u�<v�������U�o�u���N-[�y����:�su[_��&�aBiۖ���T�>{��������l�����|���ݞ���}�睛��Ƙd��4�8���W�s؍��k���|>�/�O�>e6��;w��?�c*�|��gt�S�9���*�M������/	�_ �Յ�m[...x�p���%u�����5�>�]�]������:��-QO[��.`]�Q��(�h�~��d������A��k3ʪ��o���]@>0.۟�4���k�P�=HR�e
�F�����d����([����&�Xr�&�&���_���<x���kpE�s9�1-U^2�U�U���1�_;bo/��9�+0���gR������Y��X��m[�������h�2}�=����̐)��i����o����>,^����#9U�c�Z��\�8<���o����w����m�K�~���\o�!�<�؈1?}�C���;8�����r���zï����j_W���<c�*�͆.���p�f��&���!G�`����7H�%K�A׶�8�������G�tL7XY�}9}���%ٗ8���� ��{x]Zvxn�����kw+la��4(��g��:i�h:Ď;�����1��Q��#6st"C�E��!�}�%���������L�b�f[��������%fk��4eq԰�g��ĎE��9��=!�(��?�I{�؝�v�� ����m[�>}:�F�g�`�1�F�:1�"�` ���H9[`l�f��X3�-�B��d�h�1l0����,^-j0J�5��ir��oY>=�,�4���~����}�EG�C����f�SBlh|�j�A�/����J&�e�/@
px�k��ڂ<? R�v�ɖ/u��7�^b\A�AME�w����,Ѯ�v-�2��A������f��g���~9ccN��9�+�l�D����%ưI��,�ܤ�0�1�brCk4Z�1ڦ���nr����bFפ GE��s�_���:�񂱞M��5�r���KU?@��<_|�>o�(6�>�l@�
��p��&Ȝ�7XSp�v�0�Ő�!(��D����φr�2+�v	�ѵ3j_�X��7��	��%F#y�g�>������'?ͪn�\�
(Lj�+�d�x�6o�s��|�����#��32W��!M$�>uGQO�"��
��hP��2a�˜�)MS��[�IZ���s8OC�Q�C�?C�>O�r�}%�
�:�d�b���IZ���d��to�|��>���|�,�z��<�ɭ#DM�(>��A�1�4M�E}��za�WEE��mOz}�z�K�fgq6I��2���uڶ�j����߼���|�?�����>{�����&s�����ͦ�+3��6t"񍯾z?~W�8la/�ce�|�FD�#�aA"���X�׉i�!�Eۚ��x핅R�EU�,3��JQ���Ij���O���اo����=�}�ݸñxј��#�m��دM#�ADݶ�4����G������u����E�/ұL����x�v�M ܾ6U�]}�0���W\_	=��k��9����Y�H}?SjS�퀚�ӅK��=� 2���y*�@���^�7��5j_��} 40��u��Q��,P���oB���P1� E�%��j�P٫22"��s|S��Yb�B�A'��5=���[Ӹ�=S5���c! A12�=���� b88ا����4vm��eܸ�*��������=��v�%ӂ��|�D�F%�U�K�K�["�.Y�Q��])Y8Ǭ,	]�z��,*Y��S�k�CQ� X�vM�58gp���}J ����M[?����b��n��;�?�=��&Fx������֍~��ۥ��eb�h�I��]��ד6\7�O������A�\S���\2 �ymZ�7�[_5�:����[���g5b1��ɡ9���Q�����7o�^{�����tE��˽�m�\_,�e6_/�U3�F��S#�]��߷}��oZ�����<�YQ�m��ں ����""��L�5��z��TkS�5�B�P�Fa6�spp���UUa����d��7��h�	;U��1[�U��&�]��U���tz��ƴ���s�D �l���=�Z�(��dw{���դI|��@z`���Ƌ�PI�{췟5�tL�8��ɳ�Ƨ��Ŝyf!�t�s�ӄ��D��	��:���*1�����CKQmϑ�#���Lc� &��o��Mz%VU�7c�����7߸����g�Y-ϒ�N,m���\�+'/��DC�$��{8�����oq��c��%��s�^�xM���.Ϙ-�S��$��yU�g�^�k�T���&}ڬ�ǿ��0�z}�����,�)���r���������#n�~��܁n�я��:��A�a�����7��Fb��	��J& ���4�b��%�EA����A4���;�dF��5��5upq�����`��uZ��"���Dv��a]�������$���+�͒��CL0Wҟ��cj��1q	p:�(�kDl���+��WOJ_o>�.��ʀ��D�����(} p��iX�ZxMר�m���AS;df�4n�2�޳W�Q�mӐK�yꮥ(
n�r��w���l��?��}���;˪�m��z��iV����xs1�F,D�R�ks��k�ߏ�⇻w����՘�T"�2WU��E����>-X��U��#"�,���V�#I�s�֭�a��a��i7����{fS�����Xh+��YFj�c�����/N߼<+�U�q�v�9Gx�04�쓼ܶC$qZ����4�t��)=���K���d:��}h%C��D��"}�Z�jV�����7g�<������әQ20eەί�>M�
27Ø��S�Q�d�lm�e	��{�Ǟ�S�ٜW_M�x�&U�&͕P-��!v�1��������'��G��O~��ݴ`,1
"I�Ӽ����v�dICi&�W^{���y��-�3r����ˋ�h&��U���;������<�.s4$�E�6��V$38��&,;H�-;���nY�qx��W����c*m�6V�Cn������َ��3~��_p~v�_o[f/��R����7��3�ԛ�f�D�C�;2��0b2��Q��!Y��� 6ptpȭ��̪��Wl6��I0b��XWR�,c"b<�j�!�b��eP��@Ҧ
C��T�#F�Ce$i+H,_���OÒ��jp�R�͘Aʰ6���6�S���ϧ��H���UZ�an�(����,i����ޭ��}�Âl��]H����9��1�M���s��}�3WV?��j]o]���~�)�g��wc�e�4*1�h�1��3k�ۨwZ��{��_�p�gf�����hL��Sj����^�MӠ>��ʲd�~��>�p6go��|���zk�x��#�:U����,�ެp�1�͈1�^��҃�ݔ\�BׯО��>㺆��k^�<wטy�V�<�����B�X�9�DljJ�2�y,�L}Ù�od�{ʪN#ik"\��DIiЈ����#��y��_9���#�ք����xd� 2�,2�5��%�cR��*���
4Kj[��� F|���[U!z�{�n�<���)~IYVW�EU�����w�Ƿ?�.�=���!?��O؄��ށ1U`�ʣw�1Ơ��YVp||��߾�뷎�Y^����?�A���31���f�7�88�KQkh�5{{{��-`0����O_	���`��㙼6-]<�����Yl����T`209yQ1�/8:�A����K)C1�9NZ[�1�2�~��F�f����g�c��g��,K�WԤ�cR��G�:^{�6��6�2G}@���K��ϓ$A��`�l$�8ź��<#/�5b�S�p�!���8���.
�ce��@�T�g�3�I�D�m�_�}�����W�����9�з̆������p.v37]wu�we?/Z�D�f.B?[I�碑е��,pրFnݼ��w���?;�</b�7���<+.���y>�WD1)�u�*6��uB��j>�z����~��G�_����S�}��_Z�;��9��yL���*2e�B�EA���w>��g%Gܺ�*��=���'�z�`j�P��{2��f��ގ���)=�|[�iD��1q���a��z� �E��)�ڦ@�x�=U%hD4�5�c�!�b^�bi�@���S{~�����Ę������׵!�������H�޸��������|�Wy�W�厧�����SX�3c뼘ͩf�"��e���2�8��r!�����im�y��_��[oP�
�6E�#H�>�׾hj_�GVV��TA<�ރ�ϷI4.�����⌣A>4�`]�S�%CUU,��KU1�3c�;��#J�6	��	�L� ���n6��c@���i6}���N�Pb��,m�+��;`V-�=m�4��u�Czw�L���8���F ���;䭷�Ҭ7|��4�ŇTt���8KQ��y�M���c���w��tmMY��Oy���V!.�J��,��&O����� ���#����QM�Z2l�0���P{�1p�����'�!�[�J[w�.��ldq��	�b	l��u`����|���5���W3�sS��i��U�Q|��/$�ug�hL�O5��O��{����(J�>9����N"q�}���Rڶ+˂�m��*xpV��hEPcqA� z;�����޽{'������~?�^�;==��i��<�L>#��W���1B�v���WF�$Z��#F�,fs||��|k3���X��\��|۷�I��C4U�%����*��]�]�qE,<a��c�^��{��o�
1�?ϓ�~(��7=Cd9���c��4�k��{���zI��&��F}[0��l^���&�9v?{�}���u� m�P�2I2v6��+\��Bf�TH$��9��R���$��,�c��;;�Ȅ�}�I�4-}FDȜŕe�X^\�֎�y2c���׷vm �P7�:��i���^�l6�(g�9#Ĉ5��o$��R��c:�^�8�,-�A���l:V�����-j��.x��"Y��Kתźl�oEl���4]ϔJ�K�~��1X1��IŚQ��|>6Mͦ	�Ͱ�@q��s7�����X���a�v��2��u����6
Yf�Ǽ��?���&�����%�M�k���Y-*���'|p�ۼr��1p��)���'����E��Nט�U��������v~���-��AŌڻ��h���m�R!��AcD#��Ohj75��B8�����j*n�IB�y�Wc���p���|
��ސ�麧����;D綝�ɑ�|�"�?;�Pb�Ȝasy�_���G�7o�8C[��O��������N��������w�<#s.�E�v!h�]�{�������㏟��~��ٟ��E#iܻw� ��?�?�P>��c�������R���q��I>:?��~���� �/��\������E���B��������ƍ�_{�;?ߗ��;NN��ƍ�z��}�}�������_�p��R88�{ĠbrUo��S���~t��òX�s�֫���u���s���G�D�z�O7�u��m�1��c?}nL�M������غ�z��������f��1P_��m��v|���lk����r�Z9]N���q"�5�ױ|��^t�v� ]��aHJ�^��	�5l\�!%�:�b�A7��Z�:v��k[T��4S=D�]���[Oȁ����{{{l6���3�,U��Q
8�]G�帬��H^�1���vKM���c-N����e�R E�M��,O��ITn�>X'���B$e� �Q�|ĊR��]�s�u	$���u��� z�w��	���kD$�����W:�ڵ��*�����t���mi�T�Q!
�W�=�x�=n��:o��O��qvvA�S�y�8�q�͛798z�7}Т|��O���gV���S�������MA�1�	���	D���TE�r2�0*D�
E�p/FM*��I)��Q�@��ԛ1�}��v��'#�&�gX�oȜܘ+ݛ�s�nM��� yW߷�^H
����7�րj�5�]S�b3�t�D�Ռ�����?���5~����������A_#OO��޸s��52�ϥ,�.��m�Vź��Z��e�H�T���_���|��;w�5 GG���%��������Ł�ϗ�$�I��O�	K�b�ң?�|_��������E��sa>`���ê�ͦ{s}e[�u�C��N���θ�+�r��23ޠ�>�O`��6\�����{pq�^�*��9�rpq�7n��­��m<�߿������߿��Yy ���9?7{'{�4M8�}*s���b������st�h���ߗ۷o�p~��G?x�Jl��[o������&ڼțu�:0b�*R�A:�����Z,�mZ.//q6�����.F888���z��7M}��Eu��l6ڶe�Zqzz:������*6�u]�V�Z����}��޴�j��}J��qΡ���r9�С�k Ä��y�f�T]Y�	��-��H9�HfӢ�uE�<��뚬�Fp0�G�3��E�,�g�u'�9��ֺ��m8n��� ��W`�"��U_}n�<�����()=��`�\ARu�b�@5�����:t��ia>�,g:�{M�]��D�#��o��2U�>@0`�M�L�R��:B�8���쒦IV2���N���l65y^��-�GĘ����C��7�u�|qH�>���:)��e�]�ڌ��QC@0.��L��օ@<1z��h�Z�XU%�YEa��B�ئgx�9��kW�hH�P�u-.�8#lV+�͚�zMD�7-�(P��@��*��Wdԝ��k��"v�h#1P��a}�V���xQ`T0y�KV-�z�Ū�����8���V
VB�$��ggm����5?����w���y��1mW��6MG״�9��l�ӧ?��<<�es�M�K�2����g3���8�.�H[7\�^p��w�N����999MծU�5>t=A�g5h)�=ڮ��"G������l�������Ӳ,�l6����u|���p��S��=��&۪]�����r�;��$]ښ�O��a=����2}l�Z�����m6���[�4��:}��|�T�b�mNOOx��o��W<�����=��������w�ʃ!{!���,�fM�̾��o�o�w'�?^���*Y�AbUZT���ܓN    IDATET�?tm�'���J�� Wu�ie�Xi��^D��5�w$�pb���ցD�x%8a>3�M��=Ʊ11ΈTs77̚�n�K�����;(Ķ��B̬�U~�l����n�cC�z1!�,����!�.j� ��<-��b\�}p�����y�ESA	������tvS�l�A��x�ez�7U�����N���6yfo��u�J��d�w�j���;�w�6y�m[h�7Z���E��f�eM����ʽPU��.+�B���W�;_����(��Vwſ���한��o�f�ݸ1��ixp||���������Kc��l6ݽ{�����NOO�\�5�+13Q�1b��ī��mT�n�,�x뭷p65Ä�&��׫x���(Hk�dbY�e��͆�O�r~~>�����:�Ŕ����S���޾)��g��1�u%�,��z��qS�X���)к�=F�>Ҵ-M���-Ӥ�k֯{q����n�~��b۔]�!b�	�5��8`zoH�5�0<����C_tS����`$1Y��a��5�-�RW��z�.��ζ�=�3�R��:V o{٦s�ި��*[L1DL��-$�kX�R�%M����#���p����� w۴ب��1U��3�;���,�łX���5��c��H:&�Ӵ.�)�j�6������pǤ�����g��M��)��W&y���i �@k��9���J�z�L-��J�U1�*M}��ܣk=?��g����|��R��s.�k���e�;ڮN�[��'�i�@����զtl"�b!�v��3��{�����3N>�9���}���;���Z��4�II�Ľ��>=y�_�Uj3���#.�c��̥-Cg��Q�˜�N�٩m��Bi�Ϝ�磌g�G'��4S��2�~��0�ͮ��kԍ7&U�Pׁ��u�<1�ܹ���G�����p��W8><B�ao��#O�HF��C����7����ˋ�VL�>е��T�C���\_���FI��Z�T$X�b�zb�eTD�Q%�kC1S�̚��D9��Β�J4)�*JĘ`����FUEĨ Q�	���V���ŒN�Һ�v��-&�L碪��r�ƺ`:�Y/�b�[G�FuAr��G�k�����R�h�4�t��D5��U�#&s���-vf6�"��"��\��3�f%q�\js�l�XjŬ�ܬ��;���K�ɨ8��1뎉�Hې�m^��q��q����v�7Y�B6��n6�ʲ�ks���b����7�g	٧]�uw��]��?�*��]��<W�$�6"#:rwӃ UUq���͹�\�&�ҋr��k����w���ZR����#...Fo��b��dL9�7Ֆ�����5ɼ2�N�=}�5�E�S6lH��_��_:��	�h�f#z�u�l6�Q�͚��s�����A#/��Tӹ�n��z�x ��(1M�:}��@H���\0k2��r��T[1�X�V���چ��X�X�8��t�2c,&�WR�)M�����B�5l�5���z�����'Ӱ��&{
��k��V��#Mo�������.��q����u8vb���4��L�"�u]ӵ5]S#�2G�;p=X	0wm_���
%*u����1X㈴ĘLq�
��i��8����₋�%��IkȺN�M�\"m[�&IF�u��S�r��[��g��k׬�K��a>K=�����Ԡ�>��Y�DB�@$������'_�����OL�5�\h�!lVAl9y���}�)Nj?������4�ҵB��@S�ԜG�rۉ�a�gg�|��߰٬x������O�tWto�����K=�-�؂:�I��ᗟӬ>�C]o�(�!y�7��#��LA�.H���yN����֚�|9�A�<�4ד)�{�� ���Sa���bI�<�ٌ�|��w���W_���^����6o��M����t1����l./8]y$*^��(���-2�yF"^���ω!��~�]����Uc�D��s�XH�D4@��QIii,�2�Ё�9�s�:^��X�V$��#U'`�%s���	䑪�m�UM�լJ��mG��/ۋ�.R��9��2�>7��Ġ��� �b{�U�:���;�մb��"�;�D�v�� �X���"�Y��Y�c]+F�j�1��m���a���F�"�=�EQ������i��sYQ,�z����ڍ*j�|]�<���_�9���e�֘�]ˋ%p�������������;�A_]ty��&hʠ��QTt��KF���IÓeI����X�ض�JFY�dY�GMI�W�%���G������<�5OUU�v5]׍�@�U�p|]yMY���8�U6oMi�i���Y���+����O�!�9��#��������M[P��<=;e�� �E��s`��:`�_"38v��A�b�^W$ld��WٶOz�4���ټ�xHYY�
�b�Tx;��I>���ϱB�z.�Ki��f�j���ҵ`���5l��?���c
=E,Q=b�X6�ߦ����H�3=XN��u�_�4�햳X�<�E�
_Hդ��(�Wk1
��X:�(�,+Fˌ�����O~�ӧOi}�f�b��LT�L,y,yQ�9*�xYg&Q]Had��������euq�/?��Y��3�g�,�5�I�~���)0��)_��>?��g|��_�o�;X̚�fɬܣ��j��_�C��/~�j�%_��m�@�`G�/"��Y��1F�&�8C�����˧���D����%��4W�A�8��2�|�!�D�"��߰<�P��9O�dY��U��!ec��~���y�� ՙv����{�n��c�_�6c�7����fX���dY/������o��ݻwy��w���;ܺu��2+J=z�f����������U���3�\�XV��lV�Xra��QCX��^���������Z??F�у���A�#��p�$1���hLMf2p��b���Q�_�W��!QP�H��QM^���9Y��ۜu�f�L��b����d�y�'K&�I.b2�JW���^ٴB0�"�)�N~��)�C�tmMYU�Z����QU3k��]�*s�͜u��1#��ط��?~}�f0ԛU�%d�r�]�|��c�Y��ږ�Q��W�f�Uf�jU����5��6���lfT�s�޽���/�l�ݻ�߻w�u Gu�LUz+f%BkĄ�D��$]�GP�\^^0��{V.5Zo�^�=UU�h�.�T�1z�>=���?�����o�4h�|�Z�z�M��=O�4�cl��vZmE��=�wB�� �nzy:AL��>��%Q���j�����jE�n�,/Y�V	��X|M`�<�7�+���2��1���ܚ
�5J�"5�u�=����!ڱ'��@4[K"�B�'�hVL��B������:�e;QJ��뼠�r2�h75�J�:b�p`ˎ�L���mQ0���勉�7��q���l��2�U�@LbOڶ��Ռ�#�����T�ٵ=�*F;Mc�j��ɖ4y��r��|�.�s��N��g?��䄳�?9�r�ĺ2u����9\��l�TC�^D�C_v�7ہ*����C>���'>C��e)����zY#d�u�1zbH�e-g��V,O��~Uc�ʉ�MK׮Yy��?��_��9G�ѐz��%EL�O�4�}
�<�F��<!��q���"��!u�5	XxLH�%F�@�,�-�� �ΧjQ��Q�1���t����3�������삾�rw��s�f��;�i1�n5���0v�߰�4M3j\��eYr���ַ�Ň~ȝ;wx������S�5'''<y��#'''<}�$IDbd^Udα��鹱�!����S��l"\��Ҵ�����s�ME����h�@HO�Q����'�*4>��:��#t�x�Z�HD4�&U���b�E�o���65��3��_�w�@V�bFUT	M��3��g�+	VEQfe���-���(������6_����w��	IA��-�K�f���]��B�AIsL�<Yn������9(ɒ�,
��84up�\��ǒi}�P_�Y���(1!�����ˈF���,��6�1�%��T�o����;u~����'����2zF��1ƫ�
	�mu�� �Ba-��E�et]Cy���z��Wcx���O?��Ǐ���P�8�A�T��\1J��tW�)?l�Tp;�wx}�����@�n:z؎�x�뇱��M�1�"�	1|�5��6��כ���r�Rt�b~I�;�M������a���6���k$�)�#^=�E�<g���J�M���\����V��CϘ��9g6�(���,Y.�����L[��:�+d�$1}V�zk�:�˔��6�Ib�D��A�4(W��q��A%bI��vQSM�Rg�������ᕛ7�_�Y��ҮVtю۩�	�����٘��,x��|����x�����!�͆��'�כ��i+��a��rA��1h20F�$]c:{d ���EAS.�fţ/�8y�����e�6�;3���C숱E	l��B!s�e��
�Ո˓UKpdF(r��j��X9g1��3L��&}3@DL�'�TS��JJ�9k�3A�@7�ov� A����JJGG�(iaF�,�e��Yb@b?���oۧx��9�g
�^~��n����fC����9oÜ;�����zF^7���a�If�u�W^�|�=n߾͍7!����>}������
>65��2��b��mq.�陼���e�q�&����1a�*��Ҳ}\z���ɶ
��t�-��ߢ��]��X	��q�$�g]�X�㚀!1���^�Q0�.��M�vE�>I>���l���׈��9�y�&��1cG�$ˠ���R�r���ɈJ u��yF�2��T�%�,f9�2cP�X�O��h�(+9�
K�}_f���l��|�N�1l��HJ�u�
E1��m!���9B�9���w�m �#��*���f�[%Rh�)�[���Kg�����7��w�����Y��k���άx�������N����������0ܼy8���g�<�mkNN������/��p���[am�6W�����s.//��`)B�� �)?ܘ�"��=�vR�C�7����ԎcwB�J��w������x�i/d_��,i�+��~ۺ��/;�=��{�{~�GR3���<�Ry�[6��V�`�6�O5�@:z4
y^��w�|V���M��-Ѥ~��& 7'C0Q�%7n�^�7nQO�<%����21��~���p�$M�V��h�5�Ѻ������,�Y�\'����C:�,
n�����Y-988�ެ҄�@�Oo�Q�$�#�{�=�~���{ұ����$�1E(-i1r����ʶ�r�?��'Sˏ���muM�u�[%�k�h�v�#OA`�2fW�$��X�HP:�P:a��G�u��k\!�'Ѡ�2wX�<��AN�Z�]�cj1�ơ:y+�u��H,t��(���Pa�$pb��A;\JBh�cRP#�}�qH3�y_̐�}^���~�+�kwG�7���u=ʑRox3�q�5e����7��{wg~懁�\����|�[��7��1��'D���3�e7�u?7m�]�B�D��XI�<�Ec�n��J���Df�\N�k����{'�="�:��ύq���e����Σ$#�:4B<6sxBj� 6��GZߑ�> �B*�I�#Ĉȝ�� �@��f�X!w�Xd�e�0E�Yr�a3�3��f1��t\� A!*]���:�}�5����.�t͊ns��| Đ�m�~���@^D���C�v[>��������:L�UU5� ���p�Х�S�3�/f][w��NC좏A�uU+մ���<��o�7��o���%��+������8���w��l��d��[�$˲dnC@Fd���h�Q!�4��Z@��4�Y�H��;�l+��lQdS$��*��>��{�W�����[,6�d�[\��{��s����������:3Ea����+��V��pe��$�*���6M�Ǫ�B)��#rt�<R�nx��>[�=���bI�?����G���`�e2�\.Y,}szk-��m���1m۲X��*�d��n���tQ�"���X�'ɓ���ٳ���/=�OS[j����%�"*>�inO�7��8��V+�QFf�$����c�Y s������{�?�'龒/��M��E�/]�D�:}�8�X.�ƚ⌣����^~�+7o��(�{�n'G4�5���ڹҝ�q��2v�PQ���y����-�w�,�K����R�J�㒋/b� >��3��T��v��Z�b4�=s��M^}�U�I�T5�Uloo�2��H�Ef�Hy*�1����-ٙVYgm :��m�7hi��[��� �!A"J֕�:E_T\��ʁ	ˣ9uh��꺽tr>�1�>t�!aRf���P!�+|�$��&֩O�Q�' ��������1:�I<Zi�*pc/v�`��v4�%t�U��6Fw�����E�c�>��
�g�&�;#$�EQ�sz�|��g{q|�kG���u��7"���+wS`$���Ʉ���hc*r��f�6@r ��>�9:����@T'	�x4�{߯��<���(ǔ�s�}��yR�Խ)�&b �،Q��I�Q��y/$"X�is
(��z�����fٴ�I�ת����K�M��p&�&t�=�x���m�#�Yg�T��x���!�5e�h��LG kM�mn�t�kޣ�f6_���Uv>�;�+�R��&9�J@ɺ�(ݣDq�����z��=)8(�(�Qh�O
o�|�4N���m��ku�g%)�b�7��v�g����y8���6�`�\n�j��R�a�VƳ
�� �ˣvw/���G�������oE��W��cV͌�?�1<�i�Q���NgGL�SƓ�
SJq��5���o1����8>>E)�1ާ���½C�^z�� O��4��S݀�<��M<M
k�|/����~�w�|MӰ���Ç��U��H�>Csr�À
��D���dZ��-"��c��e��e�x�����I(���ւ�&�Ef*xT�γQ&j�)>�B�&�:}�_�w��g`�g����*?EP�����Ũ1Z�)ѡ�Q84���*��U��u��	%,������� �#C�u=�t��&E>��[(�͕K/s��_���i�@�\���V�d-[eƃ�Q��'(}�>к���Ӵ�n	��V���r�EE^��$��'�a�jE�F��<�,6h2Q��튑��Tx�Ȳ��Qň���k�����OJ����]v������������#��=Gh�dh�O�=��l��K/p��7(��x�-��'ӆ��.��㼦�9:�,��� �
r��!U�nF�d��	8:�E ����ۼ~��ϗ^�1�VGp`u�!J�b�fg?���},�cE�� 0�.����%�	�Z,G�n
13��$lN���.�$	��1�����R"T�l^;�B��0�D����9�=�E)��!�t��Xaӱ]G<��iC�,�Z�3KE�6�M�~�a&�5m� �-�uEU�(��_���{ h�(�	�̡E�#}(pz�b:ً �$X����h�K��B8�+\]Q-��nUL9��<\���1h(��rdg]&J�>Z��fvtS��f��"���,�K�0:��y$�Fk���A��W��9�w=H.�H)Q�vx�����������c�AE
��cg��\W`��|ۯ��1d���sWW� �#m��s�(�ƪX���=H��#t�_�����t�������ޭy�!�u0�w bj��߭�Xkh3EU�m�〻@�n���
���g^��V>�˗������,����QZK�����/�M3k��f.�,��[���X���~[^{�TGs�:Q&[��G =�/^00R����]�ܹ�������l�����[oq��-����s����}�:y\GG3._�L��ܹs��x�o��o������1��ǜ��Fo�5�D�>�mvAaRl?������3Q��%�q�<�x��ώ�������A��/y�q�$ �g͆)���Ǒ�i��p�N$����˼��>���~��l��tL����nT�%�h¨�H��]���Q$ت!�    IDAT���ZK�t�g,΋&�s�
�����cn����I�$(��	�������C������w���s�Έw�����M�v\'7�g�$�j�(��4�(��mFcW�&�#U�f�e?�lΡ��t��j"1=�N/�E})���9�Ʉ�,��f(5�����⠦*ߴ�TŞ@�s�b,�E�&�u5M�hh�S�ȳ2�.���G�{��K��c��9�u����1%�^kF�6��!���v^��6� h��^�0�D�[���B����c!C�{T3�H}��#s�og���^i��A�1�����k͙�cHAm�ޟ��M_�Sy<�;�:Q�E1>�Q޸����sM���.�����m	N�:C�eUD��kc���7�o<J"�w�d�e$�v��܋�8�*ˊpp|�����w
�G �������?�C�]��޼Y��� �k��R��cVr�pV�>��5�����.�"G#4Պ�Ǐ����������Xr,QH#��R���n:����)z�"rC�B�*|�=o$i�����t�J���l
��0:8l�A��c�{��QA�<��8h�Fbi��l������,[�xz�*����rU�ZF�͛7��sz:��dƅ��Oڻ���uǁ�vc�w��^p.��<�êm�yG���?�����!��LS9J�H���ˎ�prr����v&ܼy������i�k[�	�CL���E�<����� ���#tabׇS8��Q�t\��6�{?c�o��yLrf<�����>�eY��|��QJWN�v`����D��<��g�1�Z6t��-�SB�ڵ����"h����ƍ�@�bQ�B��Oiac����u�u������i\gl�G0�5=�xPg�ADȳ���E�����Qx\��u:��Е�F]>m#�/�QVG�<4�9B8+~�;�f�A*���,������"Q= �MA�������ߪ;��<�FY��:��˝t��$f�b1�CY���F���mQ�>q͆�2+#�,�."�u�w��Y�ʺk�#73�U2B�m�Z�"�����o���j9�EaQ"���m���ҕ�!�6C@+����޵�Z���K�$�E�G�j�/!:h�1�`D�&`\��YU.\����;w�0��1�0�y��1"���1���K$�:����������'�'�y�7����aLy�/ے��CO�i���Mj=_�[�B���Ң:�H�{�����s�>R
$�u�Dzr������.z�7�{�5i}���{�|>����u�L��P!`MI�QAp��l	jF�j�Ν:�<~����ׂ��3.�paY���`�ym��\���s^ʳ�~wi-�c�����e���)M2.^��d2��e��:FZ��!�����f\F3���� &C�"+�vDլhR�����I�����>[�-�Zk泓/|�Cg9��ZF��ɄK�.���)B���w������D~ga��$�`�eU5� l��q��M�]��x<a:��X,9::���������+ ��M�^���3PQ4f��<���Ǒ�qڲ�k�ީ )5��1�'���(���҈�B'���X|P��<%����FcTWr���+�Gi�o�t����Q�%η��b�Z|PH��wxӤ1K �.E��&�4!X�b�������L��@b��&�,�z]�s:�E�.j9�?e�"�v8w�E����z݂5����G먣���UyL�g�}�I��EiqU̈�m��AME����V��Ѹ�W�9�ۣ�3�#�[��w^x�;��*S��sJ렻�k:r+
��'���{�6Mӟ��Ǐ{��h4:3�����t:�,�� \��q��3@+=\=PROO�~�J�{I�A�.���K��	`(�YeY��ks�9�=˪�"�@�QJ�R%�D>�ha]������'���&�,��$��v�������>�d�A9������~x�ӓ9[�����Q�)G6��E�ꆦ�c�$z���wTZ�z�ꊐ�wݤ"=Y��l(O�"���2��ֺײL �L�4��	=�{>�s������^�ҥKL&��S7B�:ڦ�Y�>�>�t���kb�m{{mjZ�ԡAw"��r��k���5�yub~�l���X�go�y����km ���ŋdY���Q/���Q�����Y�ك���O ̘��vQ�ƹ��Zr��n�x������3�{~kh[χw�X�8::���CNO�q.tѯQ&��:��d�h�Y�#%��E�b�61���T�[�4�o%��p(/��^TҴ�V�d�H�Ġ�{A;���(c��|���V�C��DmE�AD)�h|z)�D;�Ĉ��:u唏Jv�p��w������N��|'����	^�(�g��A�V���V.x	�uo&j�k��@�j� �R38F%�{q1L�<*"U!T�~QJ�6fuナ\� ��AwaU �e��Z�R!�(o��D�;g���5�5���7�m�Ci�^���~,"�d��cT�#c�_TҾ$J��.���D����+�>��ݰ���p73jn0�AS*��.�b�\�΍�e�|���I��h�?$�D�;���ӓ������dIѮaĦ���q�@�{�8�É,�8�ӳD`��ϥ�0�Coq��U^c�!S�p��'-|�&���`C��� D�D��mt6Fk������H]��{;���(�mmAS�hcQ6G)��9Y�DӇ��w'��gr����y�g�)�ϸ�O�cl3
� +��5�c��tM]S�Z��>����6#�
�wH먛��ZRU9M�p��iA	YQ��w��tBF���
��h���D�6��	"���f�yk8&���:cl����(Pb�nR�T��g�\��ߟ�'���kU��7�=/��uv���F#�˚{��������x����rA�BuC��y�Q摧�"�Q�b������x\�}������4.���*���.�j)�̓+�U�#�#"!��˃3�6�B������Ҳ����T��SA\�ֵGG{˽�����RY�}���De�5~���Yf-#�m0bt�G^S*t���8��ʊ�hU(��X�j��)�&JFi�%'�$=�L����z�u�M�h%:+�P�X<+�m;�����E0
e�Z�VDƙ!H U)%�U�P"�(gă2h���H�2�J��A�ZKP��֡PblP%�5�eZk/F0FBQ0� ^,J�,ӡm�>��Z���Ѫ��ӣ��2V�8����Ց����Z[?�,܍�dr�v��}�Mu���Fo�컂:2YvA!c"�[3�6�\p�ek:��Gwh��o�@�4<~���>ƌ�q���0Ĩ�V�>���9�ٌ�ju�T~a8mxF�睴��lP���P�~pm����I��a��a$q��F16�_�K�mʒ������OZ��l�D�(��f$@G~L/S�����M�w���{����d��$[����f��ݝ��&v�(�y^c2�9��}�ш�h�<� ��{�6���Kkr�9�{Q1kL�oK�hkk��ׯ������#<xR��0x��������-�|�2�Q��|�ֆ�V������=:�{��p^��+{>��3M���%��-t�R���u�z�g���I��'������m&*���>^�o��;o�����!��
�'�:[W��6��&F)3Ma.\�!/3&[1[���y�_�4.��yh�Z{�B+�.�������v����+���b�ֈ4���MF;�V�΍��b]v�4�,���R�UVm��.��x5*���3����o���_��Q����O�(�~�w~'�����z���۷��۷�J��}�������t��6f��R�c�ƹ�Nm�k��f`�UJ����{�L0�k� w�X�TN�h�>�,�*����*��\#�l�:d@�dNkk�C�Pʪ�����D9���s6h��Z���8��1GΙ\i��֫;T�+��*��Q=��Tv$Y�a0fi�ʴ
�m_���AV%e����t��r)�nݺ%���8��Ng�ڪ9Ɋq�> �Qd���Ն�ka�X�e{{{����������wI�(�F��szz���J)f�Y�oW��x|��ؒ,�đ�`f(�.�O�g"��?M6��w�Xd��3�9�ߔ~;����6
9λ?�`/�ֺKu@���Q�1ژNGS�N���}�o��_W4�Q�Sc3��N2�����۟Rv�q6/�F�	�������g?�R��|Ч�O�*;����"`C�+��˶��ӊ<˹|�ba�Px����b�xd���ĭ�H�{)6gw��l;�T���k��
5��Q��싷D�I4X��"�T�2�s��Ms��x|����ŋH�O���$SJ��|��z<���ϕ+W����㣏�����hm�K���!f�(W�5ň�t�h4�����x�R��|�jYc����\�x���s�}ur|��T�Tm+�r~$J���EU��AB0^���ki���Z{�6M�hT��f��*��F���fbmc��Bp&��[���=���mk�x��znL���҅������ (
;�sY6��۳���ܵE]x_Ε�lQd�z��������ʭ�n�ɤ�>�����7.2�im������ڋo��}���X?��P���M��,�q�X\�U0�h�[��º���(-
_�F�bE1c\��s����H���Y�H�@��X�\ �i��~fA+������ked$^��z�DNuΞ�m�>
5��⼘V�4�B��ʚQ�C}\Uvvv�yؒ�upppr��α������p#��TL����0S� ̛Z�(T���;��{���_����QJz�w����ۿ�ۏ�.��o�b\������-�7�#����"3�l�o�V�u��+˲�%�#�u��UJQ�%�ժo�^�6=����CUU�C��]�Uz^�^� ��� �
+��<Ŵ�a��@Z�=��E��(h۶��=L��57'�=��x�5Z"6U��^��%���15J�v��Uk�8����F����f�~Y�(�δ�Icዖ�I��kK��g|��f�=e2��)�4� ����	tc� 7e���Q\�ckk�+W�2�-K	䅉�]%�/E�Z�p���^<�|��ޅ�4����qɲ]��~�yE����bу�ƹ56�<�_���ñ�RcQX:�#�����m-��˿��_������}�փ��gJ�G��:g��*>��ӣWؾfI�u�f�b{w��w�f�4��X�������ϊsǺ�?Q/"�0F$�#1p�6���~Y��}=+���:�_����ܴ�j�Y]�MK|��y9͛OK����,��y�h ��^�\�l�e9�aݖ1uu�	����Ɍ%���;�$x�ݽmnܼ����'�����&��"0�n�H�R�՝͉�c,Yf���t�r��������a6�ك�G,���nX>>���cw�?�^�tq�T�#4{2s�}\�֞�.���i''ƴ�͛�	ʨ�6�������o-���\X�.��_�z����)��śo�)Wo�R@�}��p��������խ[�$��?�?���۷��q[����i�[�n��&��81��G�p�_v��|{�j�]��6׏.�ӫ�h�ԓ�AƩ���q+���������cK/n���T`��v�%;ń-�VK���YQ�e�L���Q�y���*7�(9����ж���8�Zoy�m�*�B�h�5tЂ<��h�WZ�v��o��.m�z�o�����t>����Z!�F{��2�����R&��y{4�O��T���O�a���_[��{�;�V�daU�em��j�7�~���P�h��L_nr!��4;/�;�NY��ʟ���j�t�Y���9���
'''����^k:�TB~�bك'�؆*	;'�2�ȟeK��	Зe�d2������O��[C~Q�����$o�sBw�ӭ>*����(3�>���u��h�B���Og��Ιυ�����|o�"�/_�j>D��Gk���}Ї������/�&t��|}���-���:��p(C��2�d���|������obm�\����w?���lxZ����Z>�w����������E��@v�.����1&>G����Z��OKe�Ά��������$���s�k�d����!t����p!"�����8�
�>�E�;ֻ��x�y�w89��M�@u��Hj�f��s��e����L&�y.Jf���?�c�֎�jI�liZ��DJ��X���/�)F�����rn"A���eL���M�����?�c� Z�Y/9�o�������7���|����}�7��称$���R�����۷o���}��Pr��n�|�p��5�����0|�ߔݺõ�b�r�ܿ~]F���|�W���C��pl ���t���N�>��ӝS٫���Ω:9��s6|��U���?s������y��ξw橺}��o����<�Gʚ�b�]���՞Blh%7Zc�A�`}�&`��k�h��k�w�F<�����-`��rN$h��$�L5}R�i8qE��QL^�P�15�NQ������������2C��tLÔ���kj���gV�ՙj�/Þ��?��he�dfY�Ot_��=�6�
8[nm�F�hm�6�茠3�����ϫ���믿��䐏��ؠ� ig�OS�𐃇�88>b{k�";�\�|��/���Ǐ1&���*�;ϔRԝZ{��t�H|��<�w^Tf�K�u�M�(�J��/�"��k�dgg�����?�0�y/8�e@�v�w�i��"g{� �/���׏�墦i<u�X,*���"����Odϊ�mF�����?�g�<ǻ���p�ĭ�4B�]���o�7�����������|7�4�`�Z�4v��4k���QOK�k�d2�{��f38==U���qۺFIl���E����p:���	�R֒�F������iZ�����~0|_YgO�ގ��O�?z��I����g�������+���%s��<�ƨ�J�C����R)2�Q�Z�c��nMQ�aUk��eC;�K?�;ϔR]A�Y��M0��)B7�L��<�{^�d2��ݻ�W6L��xs�J�F���1G_��tނ�,��������%����Z�96���4�*��E�X������|�/���������گr��>����U�B�3���̎�m�v���1<~t�������`w�W.�@fe]l�w�OM)n�Ϳ���i`o�vFg��YG���d{o��f����~�G���9M�8�ɰy�V�K�>��ݻ��ҋ\�V���u7��d�b��,+O𚂍9dy�Y ~��=o�w����ڜS�c�,J۴0P*n{8o?������4�V+NNN��&���cҧ]�γ���
���CB�y���h΂�$ӚR�%�{i۶�C���'�h1����g(,J.�c�Wa�X�Z��d��3<R{q6�^�ܮ����m���৛��ʾ4{�]�������r��ҏ�׳�LByn��+q���J�]2�c�$�`:O{_Q� k�6�Ki�a�5�!P��_.����V+����,y��^���i�i�3�жѻLಪ�/�����yD��'"}S��z�I�y-ݯ3i�n<E'%�)�����C2��6.\�7�7�������_��`�b9c����g��aC�����֭��؞��۾��9��Q�m싊���o���y�/����`��˛�g�=sJAQ�i}�,snܸ��70�PN�������o�X,��#�#vDц�4e��ʐ����#>��C2{�����or��/]�i�?�׊�d�	J������m��l)�5���ߟi���cꪔ։��e���\9
|^��M��2<uS�C��4��?+�w68��{�ɘ��^P�X�����Ƭ���Y��3�ǣޑv��Ѩ�(��Չ��RH7g��hC�EY���2�2U(�[�!s^�9���+�[b�&n��xG�2[��X	�f�F��|�t�Z)b;�4 7���;�"d�҃�"�	��7�<ͳ�\7ӥ�{m��)�ato�In�tC,�3&�oP)�w	FiA�.    IDATӾ7�߰(%�y7���h;oR�=+���Y��t�S4�y�3��m�c)�O)E7���Y���7n����_g:���ጻ����!YfP��9(-X�	ƠuL�<z��*ߡ^�ܿ�|���'�FP%����;�?��7ql����.��9[�z#}��4M�`y��5~����|�"Vû?>������?��>~�̒)�hd�@��Sa�Ay�.�?�����-9x|��l�h4�,&�W(,Zٙ����7�=o�����p���,����9t��Na����f��y�O��l:��U��c�ٌ�ry&��|<��[k��f}�.�S�EQ�Y;����4���c�t�I<�bKw��'`��G~�24MMTԳ4�w>2A�w����n��~�\�W�sjO��۷o�����!�V��^�6<ԙ�����iM�7Z��(5&�Ch�p�I`( �1*6D�]oǓ���dO{�Ҥ��KO�WaO�o��H�Q�}��[)�Wo��䱹X�m�^O0���,��Eq���ާ�__��霡�7k�N��p.6d�&��O��^Rᣏ>���j5�YΩ��Ѹ@���V�k5�讗��Ǉ8_��c��X�>�YE���t�U��F����ؤ(el�A*�\t�3 �<�T��F��OkM[�k����h�[o�xp�.o��gܿ�6����N,�<뜥��tJ2Z�@k�.62OQ�?�˟��g<f�#��P�<'�3$(��i��r�i87�\W���6���������O�<?3G� @KmS=1ߧ�|E`������t�S6g<#"=��yl�����ޡX� �@p�.�F��J89>\GJ�fT���m��bբ�� �
�VC%
Oӈ4M�
�[�L�Q���vF�90����)����,ٹ�Q�])k3/.��Pg�}O���J�Q!`�����d�ė�b�C/FDX���Drvayz���8�D�6��":	�=�Xy����XP�0�����0�;�,�g�����E)�{iC�/Ҟ�>P6��I�NW�ŧZ&"]�óܸ4�b���µt�)�lmm���͏~�#�̀��oO�u�B�Z�� �Y����s���|q�X�W��bww�</�>�is*g�>��,�"{���oq�ٟz�r7>7�8&�	����~������7?�G�<E�S������kY�jl&��S�(�w���ȩ�#���ׯ_�������cr���?�B���3�u���
�}
�S)c��E�R}TjHU9�c�4J�$@5�N�N��-e�Ζ$��|>�[�����9�a�#�L�,���<U�9���L��s��i�_k���.�l����YUUvMJk����s����s����S���i����Yn�	M���Z��nf�}��>z�b���g��}������~5b�߹2��������B����4���]�[�Xm0��j�kO#^<"�F���-1�:*yV���U�j)�:�������kc����<�ŝ��j�a� .�u ��􈭭-��'��R�5Vk��8�Hal���m��2�=H�w����
)LqH^e�Mn���� ��7����0�>�i=�d!�I}}4J�j�r ��/h��>��� �8�ٚ쓛-�Q��&4\���G�,���;�2C9�?~Ŀ{��</��?<,
l�i١�u���/��ͪ�����7�������]>:XB�^�ԒǇf^�ƉB5�,���	�v�-7a��<^=�n�r˪
 ��Ni���g_�O�JYT�G.��R�j>CG�ۓ4C��j��j��
5���|�Ο>)�n����F��j9��Rж5Yn�ti�w����?�x睿���nG<<<��m#���B>�3���sC�t4M���1���$m<��=3(�S�Q��ի�2�@�C���D�z�jǣW-A��8��*�0�,���S�4ԋ9�լ�m
<��&�B�0
�P�סu���in��]�������傼(#y�	�B�`	m�$p��un\����.{��\��C�@�\��T�GǏx��!����v��Op��K�0s-��2�C�U%˓%EQ����o�̅+���,�(Ǹ���vI�.��ӓ����]��>��	�r�xOfGhM�'�ھ�Py=�k���<!�E��W>�Q����1��h�s�����a:����@�E��<��IAr(�����@C���-J �Q�f�aœ�����Jk��y��"u���N���Zw����P����xoG�z����Bi�l�������WK7�������O���~��\���o���=�2f>.���j��^cj����5֢۞ �4C~�Zb��^P	��k3D�D�C���Z�x�}�6ӌ�s���\��e�G6�|J�*�,�X,,f�u]������"ҡ� n� V���(Sqq={��@Қ�xn���m3f�%J��Ձ�N���E^���SLE����Ÿkf�Tt(��歚Nݿm[=���½{�x��8<<�Q�=��hU�V�cMp:>'*�d*�x|h#�V!v�t��QT֩<?;�ƒ�%Fg�ҢM��nɣ�����)A��Ϣ��o3M)�	����߽�|�[����V@��ҁb�T��}�"	���"Q�B�M4����{���(���X,���u��^`o\P��`��9_�3�/m�B\�t�Wn\���q+�ݿÝ��`��j(EfKP��n"�����y���y������&�g�2�h%T�mUst��;����ŝ�����4%(KnZ%,]|V��x'x߲XԼ�����_����Wٿ��YD7�x�i��+����f4.�t���O���(�5�J��by��<�j��ß��ݼW�"��66i=ß�s����q�7�g���3���y�X�VH:x%X��"�y�T"�{�ӗY�ʾT;�����w�w�R��j]XV�f�ng6�&
�ɛ8I�c����'GqR�s�s)-���#�=@���
��k#�>����,A{�Ɉ\�OJ����ސ��Ep�6�DHN���x�ŋ�����?11}��������*bH�D%@�z.�����M��"�i�g4)Ȋ��������A+E�6<>����9	
c�و<O|��H=��aZ�1���,�Պ���>"�:�y�5
�"�4�AO^(l�vEۮ�"A;R"@z�;x�"�@��1�"(�r���+��w9\T,jG��,��UZE�a���go�c�a�~W<�bXձ��6�ۮH�K�� �G�b�QxeQ0Oy�k/�5E� �N����� l��2���ɚ�y����y�+��/�2�ܼ��*��>b1?��g���2d��ʫ����_�����^���S�?z�S-�q���-m�	W.]�՗�ί�����.��۱���)Ah]C>�c4Q�w���^fz�
[��x�wx��~��f��[�LV /�g/�t��|�;|���foo����и��ű� �5�0��^�0#���������;�NN��PZ�q�i7u�L�9�)���?�o��͹<�p�t�a�es�ߔ��<��-��=�:쬳XA���������n�h��X�쩒���X���$��|��Ai��u���kk�1z�m�A�A	��Q8g�u�IWu�G)Aa	�j��;#��^��<'���R�^a�Le>˞
��0���,)ҧ�ꏡ(
F���詀��MЗ������C�}q�TmC�^^��#��.b
��e����%`��Y�,�Ե4��j���Y��������������hM�+DJ�(�#]a��6Ɠ���5M��iWx�PZ�Fx�vh1���6*�"|�Y�"���`���~�%����:�V��h�Q�z[(�� �Ƣ�b�d4B�15�X�Ed5>�h��]L�J�Պڭ�m�����h[b�a�j����7��˯p���fww7F�f�UL�F :-��ŗ`"IX{0?)�6�[��ï�������������d>;��Š�k�< ��1Fs�����7��.�v�l9c��Ĭ:F���-uAqq����_�W�W���+��&�^@p��r/�����/��7v(&Q�6*�����T�C���8/�G�ܸ����	W/\fog	-u�6��и�v9��
�������gS��0.�@��f'BL�~��Ր��C����E�Σ�9����S@�y������y�o�3�u��:�"H�v�!�J@9	�&�p��͚�~����?����o�=��1Yݢ�Jk�k�2c�dJ�1F4�#)��#h!�yDp.����ćF��Ak,��`i��0x�o�x � 7�~'��>�ڞ�4]c	Lӿ�ņ�J��$�Vp���{�r���Çgdl6���P�ŚD����F�I�9��9Z�Bق����Q�y���Kr���LIKp��b^��(���2��5���D�5dV����P�U{���J)���L�#7��ޔk�.q��.���|M�V�m�-YG��#�炀����F��4��1P�kF�l��/q�i�Nv8||����U�����,Fi�����(�mc�⪉�������zE�j2cMs�<��CPh�c���=Ⅻ�^����J��y��&���Q)eh�Z#�}����X�<�(A�`�G�B���/���OQ�(�c����X���~�ݷ��|4���m(Fc�|L�!
��,˹v�*�x������%���K<ZTg���%�k9��|7���)�\�V���3޽JZ�|t�YՐ#P9�5��������^~�reP
��������G�G�mC����/39�Ɉݝ�}��Qd}��J��ɊŲ��ʀB�|����v�{Ӝ�Y��>;�^�y�\<�T?�ZO��͵j��u����ӂɩ\��UW葧�� J�	��ҥ����9���SA�t��
?E�Z+'(U�km�3�kl0J�lv&2`�A$j�:�����K�$Yz����9����wuW?���ְ���%��� �=;o	A� -�!�` pe�2�YX^p�	�m@/J�!��GwOO�����Uu�73#��yq�䍛uoU7��d��
�73#22"�9�������-�@���:�Օ�1�Cx���Y��QL�~Ƹ~��#-k1N��_�����Q�ũ��l�<����9�#��:��?�������C'����#b�H�KPK9�������X.��)�E�`)�
c�we��'%��s��rs��Qb����I��.m�0�l0T�0��h4�Kk˽�q�˗np��y��g����7�d���_]�J>����EL����I�=J}qcs��|�p�ڳ)�8D��'�]���gOJY���ރF�g�J�i�PVfU�j�X�P�:b0����U�=��te��J��bZ����3 �g�N_�S�&0m��\�h4��2�3JYV�;����7���J�RVc�rD�=��PE1��¸������3����u~�������rI�l�}�}>���N7א���a
�_�t�+W�����-`�\����K�ˇL���/�����+��ʷ��[��)�o}��������98�vc���/"EQ�������y���v��8��mv/^e����]���"�)}�qWb���K�
ﮏ�}w���y��������z�����ѩ�ߕ�;zdH6W�"bQUU4�Z5z4n(ԟ����s�ν؛��Z/��}a��3co�m�s�)�(��9��t��J���w6 5mk��E�D�K���H�1�`�0,+$*N�%��@�Ā3��Y�!>d��Ͼ���\w�㶼�<��C�GGG�t�<�f0�߶���&�Riׁ��`��m���FM�%�sn�s�����J�}�l�Mݲ���ݻ{�
;��xV�.]۬�	+Ч��iq ���KBlq�d<�Q8<�5���8�M�֭�%.^��d���&��$�C�E�jf��>�I��"R�c&�{�
�VL6�lo]F�"QY��n�,����QU
SR�I���RU����!��h �jD
���\��<>�2������������Z�����M|���>{g��I"Q��;��u��-��Q��5X�OKA�C%�
'a����}��6��!"W�6D"1%�p��3�ʯ�:������K������O�џ�	��G?���vl2�.js��5�?�W�^��SOq��5F�1bK6����"BԂKW��ܳ/R�D,�ٌ�{w���ko������-���&��5%�bI]�4���hƅ;�%˺�	��{b:���~�+s�	� ���t�����C��}����,JN��o�m�����$2%͓�gy���Ĭ�`�QUkQ���drG���>�_��{,�Ȅ8�ʌ���ZS8k�%���%%�cde��5{����a�M�W��6���H�'�/UU�,ND�ˎ�Xc1ƥRf��x��]ξ�o?���[�,�lv�}ܶ����{�eh7��N���b��&r���K@&�ʔm�dB����q��1���|�!��S�o��{�S�<�g�c��˲�{���3k�K99��ǄV�u���>]�[#�2�&4M�F��h�h@KP�2������4��A����ѷ�2����D\$i�<�2�UИ��'��Պqs"��1eK�l_�m�$��u�\�b�2`d@�J�6�\
�p��*B<Fc�].8����s��]��T�b:	 ��sR:>��>9-9H�YV�)kN��m<��X�X�<�����&��J'k(�u]��[�˖��&/\��g^d���t:���f�C���Sn߾���>�����m�CX[P�wo}ć����6�x�%�ַ�|�
���8%�u��α�{���m���dv��{��[?{��{��G�!˦A���1��n�ܾ=���?z�g�~�ͭ��r���f�(+�i��|U�	���?uz{l]߼9{��b�:&�,�^�`���w���=�x�DE>���:8@0ƢQ��v��_E�R%�D���Ύ���~�'�Ϩ����vt8�gM�=k�;�^i0Rc�#"FL)��J͔eM�4+M�b�|DGa�Ŵ�8����""�(J.^�e2���ܺu���^R/	D���c�i�"��!�&su��pѯ�����2�=a��\[��s���#�1������ں�p������:)+&Q����س���0'GN'z�y�
���������h�ӕV�@J����ضH(\b����рyL�\)��M��[�a8�����'+��n��8�1 ��;e�Z8V�C
/+Mwo��Ꚏ*�7K��1�+�i*�7M�~�l6��n�[�PR/�(�sx�4MK���ǶAU���D�+���9��7_��o0�G�.��쀪�N��|�g�í�e*�ý�/�u��da����Cvv�S��b��(-�G<x�[4�&��WQ-9>�r���y�m�}�����K	56շ���CmQ0�����9�� �:A}��e�6*M�1�g�)lnm�s%��m��j�]��E�@?����@z��j��E�z�iA��2ٚ�c
��A5�i<�3�^��_�����[�mˤ2�P�Ĕ�g$`բ&�1P����s|��k׮��������p<_b���X�h��b�p��.�i����7�:GӇ��nP7��2�r�bI�m�lǷs>����xT[�-U��	��<9RSũ1W$�D/�G��yj�����y��7����!���:����>˷n�����~�мȄ����,%��x�����}k�rs|h՘I�X�{�������O��l��v.�{8(Km��
�p��ڐqU�Y�$�u֡eI)d��]�<�U��2Q��M�\��G+�(J��91����
��|�lv���>�	�BI�xM{��D��:\�J��9]�w2��t�MӜ���癥˝438ι�d��Nw�0s�n���}��u&��?���w>��x��d��Y���b[\QUɠ5qUFsU8Z��)��{̎7G���e6�i�}�w�������Z���Cb�b��Sɶ���~�V�6��9�H)�v ��K��=    IDAT�󂢌-U%XI�/�7��t������;<|pH�R�$6Ɉ�J7}:���Jr��pq4>�w���$�����`�h4�(�����Ո�0��T�w~���D۶�*�*��?{t�\��loo2W��o�펊���/��4�n��0;f6;b1��6e:we���;I��E�^(�c��=	��i�R�PI�
Ԓ3�U�O�7�O$QM�1��TU���:��,.��Р0�D�cQ�?#VI K��t��3��z�J
=��!�HE.	��ǧ�j�d�N���X�Q<�E4�8�H�^Z�5�%kEmm�$��j����t���ھ.�_1���]_4��4��c�z������L�X��;�(0��e2�P���EY��D�BB�T�W�bF�������k�w�F0��11��Q�D���F�Z�4���UgQ$�rY�U�ӦiXV	��m �S�0�k;R�i��׾��?���O:}���aDR1�ު(w³(�b�Aۦ�;;;lmmqtt�b�X�Ķm;�x����\E�{��Y?��V�
�e&�_�h�#��We��t~}��1�����1�q:��y���E7����ĉ��9�>������m�z�`9;bw{�A����s����{g���;;h���뀿[M^Ʉ|�Y���xc�y�Z�A���Bo`���r�<-���$c0�uK��>;:���!���L�3�`�vL4�95!�Y[1)�0� Q�<�xz��9�-0Q-�VT� ���E\ǔ��I�o�G~ͷ'���S�J6|��U)DS�w�UG���,t�p�V��(	�&�G�g"_�nO@�k�K�jQ,F\yS���ֽd��<݌@V��dEJt�
bH�;yIo
�����&�Fl�RFULt��$�M獧���g�@��1QM��Jʚκ�cҼ��P�t�"���,M���,@S���M ���q���5ޮGU��Ԭ�^`92c�5��n~����������"�ۧ���{#Glr���QըF뽯���u�ʐ��Ȣ��E�	��_��{���l��h��kj��%�+�����v,e-�25�%�cM��5���q�Ĺ%m�2_$/�A5�m��a8�
A5p�������H
��h�Ƞ�VN�3Eߟt�d�Y3`i����]nܸ����*���F���E~����_~���x�^Ɯ�M��h֍���5?i�R=�˸��g���iO�%j0�+�6��xk~ĝ�c2�ę��#�z��E�.��{{ܽ}���}Ignӵm�l��9W��k��m0�~N�6m۲\���6)S]�ǇH��mX֋�6��i��b!�[�,ʑ�M�H�,��(�/+�(!%�4
�8*�E:%z��6�3��$4���,yf�������мc<M޳�kڦI��8��J�� �rzA#^#�J���q�"Z̟�v�IF}��tL�t�F��
���n��u��Xm�+!�)�!/Z,��t/�x��K<��M�Ĕ++練}W��9���Mn�!��_����
�I�e@L�J$6(.�-&� �&�W:��*B�#`L��e��"]Vsx����[N���n��[�������ϓ���s]β��gK����)���0�/�1X�Iy�Q���c�Z��n��E�|�>f{|��L#VU��Ԃ4U�/A*��t2J�Z�B0�	>�"cbǊxr�+�sFՈ�p���)ꔭ�Lg�<����w���/pt����{��ݻO��:��N�/�Ϭ^�~�Y�,��B飣���N2�����ѩ��l���������s������ڧ~�3y"�p8d�X��˙A:I��x�ܕ��E��ΘNۗ�K!�\*ki5�8>`~t�C[a)� �6+0mM��ђ��Bʮ�!���٧��������LA�����m�jB\"&�
�u��䶟����Ҙ�#c�M���q�BL���R�T��K����4�,��X�5.U=),QS�L2>VK
�8Q:�����
N��Oq��º�C3�C����FYU����X��;�I��<�:�b�ˠ����}��
	jL-&`5M���N�������8�>�n��A�²��&+�&�E�H�`<I���\�P�3�M,�1մ��k�twh'l�E�I�ӗڸB��x���S�IxS�t����(�2(v�7џofVK�'KD냾�����Y������������r��Fl��}F����''�ϸn������*Re��,�ъ��x�4"̌m� �ۋ/BVߗ�c�'0}����j�O6�F�xYSv���F�R�
c|xR6�����e�hV����;;;���k��|�����&�	ՠd>����z�rѰ�l�8�V�&`U�,��Z,+�g�a>�����b���J��[���j 'U�4�c�`-gg@����,DO��;k@�"��~[�5��1i�������&�D�3����%�8l!�o!�
�@�HL��F�h1��L�E�4I�^�hh�TǖΔW*��^*�
E�S�$��İ�N����Θ��Y���ghi�b���,�N.�ze(��I�H,F�Nq�{�*u8Xy��{?�IY�Ic�!z��4�jK@ X�8���s1�b
�kH��D�X��[@�O��c�u�}&��l�2}��AC�}]���L{��r
�����jNd�;��a�3U�0E2�&U��@$1	$ÞH4i�ŷ�U�FD�">���b,���B��+�gH���;�]�ݑ���%1��0�C����I�Zs��Op��Aߺ�V��y��o��|ǘ��ׯǩk���~\����i�q���y��ַx*�3j���j�Xc�a�%\d��b���e�B�sA�tzE'�N��G�APO�����?��
VI�&�
]�\��c�cc#�lU���[o��o���\�t)�������������Y��(���T�N��*v<|�p�Y8Y�z�W���;d��3v�w�W�9�������'2g��Hh��h���Q����t��<��}���_����=�ɞ@m�]b�Jg!�2݌PR�Lh �� &`b��M�8am7%��b�w�o�k���_R�S
o�t��$�� I�
�J�4D�D�'��N�f|X"�슧��$���O�7&%�k*����Đ,[\WMG5%�� ��R=\���c�`�&�!�im���&��ݦ'T�vá!�F���\������`pj1e2ê�Đ�N�Q�m�����y��;o���k����U4'a���8�l]�Q���5�+�䟙A����S߰ޘ�?v�tw]��d�1�99^%%Y3�W�I [$+��eW
7{T��>g5,��[,�.�����9Gi�� �l� /�'����xw�+C,>+Ě�=u��`�ց�Y���y��B��\g,}g�c���+���`DUV8c�1VC�qv�"�p�h���wŪ�K���Q;�]�:��=E%���Ah�8#���t��-���v��y��:�`���dBU*GG3�ۻ�|�����Y,�Õ�i8��/r��e�����Ν;ܿ�}ˠ([f��t��2C���2c�����fh��B�n������g ��������=�!�b�l+�{�;�}ј>��][�+TU��]�P����6��EA-��o�-�2o�nM��dԢ>U��@��r5=�F��d�L
u:��&9ƈ+:v%�41R��#�׮�+�����	��~��VU�eC�6����/`�`]�(�.I:B��[ �`c��h}
����m��ʤ}5��>�QbL�/�`�+Ř&OԆб����;�I��bt���A'��+�>�?�yzb����*���#�rw������YgwO�k<m��+2�H�L�QQb�ћ�`�bR}��'�I���+ �IV+10'�;�poDc���KC�I��;O�|�������y5�巜��b��cy���g�}r<���g�_;+BsV�(��o}ΥJ5!x�5��c��	M�����7����:Ř�&�2)�������S���l��v.�����`&1�E0�F5�^�7���Ƙ�~���0��T3�<Bh}b%�j'�� t���hs��9f4����n�������&}t����՗~���[�xq����|���{�{ꕯ��dbT�|��+�NUW>Wg��+�]�;:���1��:r��#�����~ˬ�j2�uα������
�>n[���xU�7g��{�U��mR��xT<1Z����)�	��XpE ���`:;��E�	��]����g�V�ڝ�'�W�0�_�Aȓ�Y�K����d���pJ��Ԩ`I7�ѐ&�2�P#fD�w�ͥ-��UI��v�%b��u��<?�k�1��u����Y�_ak�E��t�DR �m�K�S���z�fxW�s���哄���bd�)7���@}�n��ۯT���-��6������^q��?IX���%v �v��4�$�r:�#���	gA�S�$�W�����L2���OK3�B�k��}���V�# �&��9,i0EEӂ1���@S3
���x��2��c��q3�2�7"C���K�_-�À-��Ō�[;4�R�kv'����fH45�)� Ô��˸�|��h�u����#��c��,��.N4�����$��˼�`��d��Ax�jk�p��.1�0��l�mB;$ĂڍY6J�~���­Ch:_)TlWkA�I�$1B�uZ�k��0� 堢�*|�Kf�}"�_�3g[٫/�Z��!�r�Hظ������]���ǝ
g$�B�S�Nk	�j
��q�H��4���E]����;\�t����������=�/�����s3�y�g����'�����v.���ى��)�߫�jEP�Jie���Z��:��F�;���3�-988�iF���!��>/�r���vvv)˂�tJ}����ի<���:�����c{{����GB�O
q�5�v,ow�����}��Y�3y^8W�;�ugc~��
f`��/g\gP�}���U�izN��az�?�cߏ=�!�I^��ʧ<���X
�)}�#�Y��[���Y�~���)���0L�9}?���HA�z
�Pز hK �k�C66��-8n����[���g,.\����|�%�ج@*�&�RT�;�`c�.�YR��;u����u�����\nQu�M=��=�/]WO���!ee�L�eX��;�0�K�zsG<s�;�Z�s/��rx��ͯ��W��
�+,�����~�[�7�~`o_��,��a�F8��J�X ����嫴m���{\�v��}����w|�W���Wee�����@#
[h1qf�x��ח���}����޸q#�m�y��"� RkJ���j	�Ɵ��q��t��2w^�	�3�p||̃���u�dr��G����?���o������.�����Y�7����ڒ�(�r�J�]FȜ���AOX�Eǯ���?p��?�K:��b�&�����	wbS��?z�EO�B�߳b8�4(<�~�-��-�b�2�z&�K�^�������|+u��3e�ѝ�~XىH*��=�V3]U��kҎN��S���i��o]�q�ϟ��ڢ#	�Y%���$��n�,V�,�Q���zl9fs��q���!���H���%֕X;���H`<��5�˲iPM����Г,�Q���%���P�����"4U�1����s�uU+X�5���Z���5��%�	��)�%A5���#�0/'�Q^�k�>%Jb���'2����_�>���l$��_�i�@-�������K����?]��ܿ9Y�w6Mr��
<>$������D,��ߥ������7�����d2����?���q|<�M��EӴeYVQ���HlU�i[��b{���e�B��f�n,74�&��H[�i)2G�RU[M��QU��VTN�T���:����ASČ�Ѫ�fs��e��px���k��s��U9fP�����N�ݻǝ;w�L&\�|y�ӛN��t�>K�;t������ߏ�v���e��������}��{���_�c��S@����ǲggl��j}���Q��S!���>}-c��O�2I�g��u��|҈����Gx���u���y��9�><���Re��>(����@��{��k���>���a�/:�%��D��/����S�K�� e�ŕ�np��5����̨�c���S�o]�JA3]2Y���_����M�B��*��O-z��uD1x�D
p�M�Z��hLY�ƭ�_�釣f��	3���@�E�Lb���'[1�k�@�!�-�Iv�j�	,j��骫��-�O�����\�u�����Z\���~��>@̥<�����=�#V�QJ�����ژ�)۵L��Q��)�[�<���/\��'���w�r6��?�F�F����g���x��F�>�H�=
?���ѧ+��e�\�sA���������E�:�u!%nȑ��*^U�*ASC:C�U�w\�L�ٳ.�RX̑+z�z2r��-<x���6��&��pLQ�)}�����u��i9��[o�|���z���:��g�2�9��Fn��C#9�7�����~bM^M�e���+�Ē��	[�uF\�7V�I��=������$�������r'ӌ����g9�kǄ���:)������}Z��^D#���]Z���Q}K[/y�͟���S�˘a�`p���ã��ܾ���87dkwL�i��-�������z�Kw��!������wߡnTO<��GZ�u#�@aS8�,u��:eoc@R&��l�O��1�_;C��5��B��s0E�+�P�T�ͤ�Wlh0aLԐ�=1Dծ�!����h��2�N��9ۍ��>�g��_�������Ҝ�ѷnY�w�y����Ǔc:�8{�����n�m�(+bT�&�o����ʵ�?�\�����H}�\��nx�޽�nw�b[��C���zUDE<Q�3eq��|��l�������_��M�֭[�+���\}�@����s( ��X�u��ߏ/����֭[���y����:��DD��?��qm�M�����j��F�eT���P��,����h��S�C�D-֔�XB�GC����������
�;W�پĻ�!����)}`��p8<�1�����H�|>˗�� �Y����ڼ�q���g���Z�h�rD�g�����w<-⪪��+�׿&�0��^*��=f)�(�~�TI��\������|�Ӯ��J�;���߫��||$�˓��'�\��˳&�_�w��67-Plʎ]},US����o�����h��k�|q¥���R�Qmy�����!�1�ł��+|����W����x�*�shU�\.�O?�?�ɏiB��
TQ">*MT�
;�nCD�g-Zv�%��Rv�*���m[�!/^d{{���ͭ{�C��� !�H*|]PT#�	�(Y�|hS�{R�$�HO;7�L&���7(˒�tʻ������^i���c_�@__j����c�ia݄߯�;�{�f�8��eM��,K~�6�ؓ��k�4�C~���L�\��'�p?�?8�z��O_ڽ�Еû�ãoq�������j��h�r����[���h�Ϭݼy�ܺu��n���op��ݹuK�_��@�y�62����U�P_���o~��͛E�M�`n޼�_}�U{�?������~n޼i�� ������z�Bw�N/\������E�p�:���������Z������GGGᥗ^
���w�<�����h���=�;1s�F�CsT�&����#�:�(�ӝiW1ã*X���\��y�7�/�گ��y���b�Ac�2/��-�����{R{�w��Px�wvFf���5g�<x�ߵ���qL�)���`���$\*g��_t��y+P�\.QMY���'��V�	����S���~���7��-�� ��#�r�9�ڱ)�I?`�Y1ۻf����2G_��2w>�
�/��ϻ�?��!��W{Xm�g����N��bwW�    IDAT4�����#�#�[�O1(6�r��(����;���䭷ޢY(UUp�+7��K�o��l����H��1}x��������oػ� �A ��5���BU�o_��Oږ��i��!��t��6b�ٚln������K/q��U�����kNk���h�����l��:L�lm]��s_g��s����ǀ�M,�I�ڳ'��W�~�:/����ܺ�Ç�<|��Tbŧm}��^�2��斫>��]x���ni���]���Z��p����e�z
�|�"O?�����)�W�v.����u��ۣ���xn6�Q�����L�b�+e��Ԉs�w6P�!L�o�����oKR0����s�)�[G
��`�;qoq���u�������9Y�	M�������^{I ^~�u��n��@���\}�+����Ķ�9޺  ��L���y� 	����tl�) �	5Ќ���rA�����a	j�_w�E#/����͛���~�e�������a�ؿ��! �H|(�O��ݺ��2ڑa�?*b�{��{�˲�"��Ht�;Ｃ�������Q�����*�(��XЗm[ԧ��"RG�V���q5	�����V�ie����{�:	�@c�唷�~���S��;���[��S��s1�#��h%�=ku��t<쭷?Zg��]}֭�ֿ���yL��1�u\^��_�X�����e��gn_{6g�>�=)@���p�դKD4yΉb���c"��H�!gN>��i&]b��~�_��3}�x@��:���{�G>z:�:�/�b�̧kc��ܹ��]�Ե�\�x��4lo�p�ZIQ9666Mvy��wU��o�5~�����+ϲ�<�ǲ�y�����������}���6�MR����Mb�)�Ոrc�_�֯����o���t�ҕUJ�e5dkk7��+��7 �@m����ä�>�|���]��$F��f1]�8^��������o�w�"|���⒢H �(
&�	���\�t�o��5~�~�?��0������>n>��>�̶]}��`�<�:�1��<+�t^;}_w��c@4U�bS�GUÊ�W�����ln�|$���უm�}�k�ݿ����n򢭎�iƣ����LhC�3�R]e�b�����=�'���?��!$���͛�$z~FK���^{�%y����֭kr��m���y/ ��Ƽ��X.2fr<��ӳ�����/����D_~�o2�V�.����`�z^/���E]U	��K��+��m�r�	UY��~$US�c$ �F�	CY��m!�h����y�^T��j��ea$V���R�S6�����Z놮D����V���6ŊB)��.RH�"Έ�a��Ęo�����b�ۑ�'������'���B�Z;zX�U�����w���p��M��},���ى͝&�u,�SU�ѫq� j�i�v�VVˢ�Nb*��M�u]�4~e2�+g@�6�L�]' bp�ć��Q�;��|�`g�2/��Uvw�y��w1����,w������u�v���s�}�m��Ϯ�;�\U�{�r�\���5�����e}[Q$ֳm�UH83b1��NF�`�;N�
ׁ�,`N,ʲ<��}�����{�o_�G�1����Ζ�@�7bp�2���FTU�tz��d�]��K�1����*��E��
cW��'"kш5��#��ćh��I�v�-���A}�hR��q��x߅�K��&����Or͞t}�lE������-"�!����bڞ������-t>	�[�3��;�N��s'>�"�����.Z�3�#�{o�.���=�ۿ��F�S�����n<��zIeGLƻ8�}H3S�7�����������3��S�uq�+*�Ұ��.��?�{̷�_|���A��k_�j0fk�����0XW�\IQ���^���*���7ٹ��r�d>�a������w��.���7�b��Ʒ�O_c:m�ؾ�׿Qp��g���}�>����C*�E�
����|�2[[[�E�1p8=��*�޽�|����vY�ZV�zHz"��L@���u]3�1�HF�ѩHD#�}z=���#��xU-*'�d�轧��GBh1&eE���`�*bPE:�m�0���~1�l>}�ҥK����O�H��������ϗ�[�������m1jcۺi6
W��Ъ��^����v����տ3�b�x��A������W����#�o���@ �������ZJU��V�TE-m��Jdo[vؚ�u^���G�~;��33�@G�)�V�h�������j�6�+�_�儉�M�)CJ��z�CE��h�X34"v�Ī�¨1�Ɏ1&��� �1��Hcw��UF�h�NJ)��F�T�7Vŕ��B�
����/��FS1B�9QI��(�b.����c�U��{�1��J�$��9KԈj"��%�?>|��;��f0(k���]1o�{�e�����"��q����UUm�����><��������$�I�[BC�Ӂ>�^��v~mXn�@c�m�aU�@V�x�z�]g�B����|���ĸĺ���>��./�E�r�h4�|��+'4џ�2HȃK�Ԝ�zM�>y�/Z�����BL!#��d�cS��XGaEY��mp�`�T<=�7]	��q&�+�D�U$U�ǈ���U�j�&��Ŋ������CK��}g,���kJ�݂��l
s�Ɣ)fU�U>3���o�"��b�w ��j��ekg�2��$@2��Z��cm�u��^��Oh�oN_������u%��h v,r��p�w���w�������T�
��&4QM��p��S1,+ں�駟fcc�b����|�������m=�G�6�2�Lx��g���a�\�\Ԉ�ˆ����~�����m��Q�>���{�R��_cwg���-�����6�����W��K�N�-'c[�-���9��o�����'��5=�ym��}4�����0�%8���m������?3��W���̋Yc��g
���ǖ�%�,Q�:���Y̗�8t�����n�_�n�AU��h4x� �/^ؖ��-�ҍ��[ΚƔ�T��Q���F5�\�/Ն�YiŗfWd1Y.mٌb#��P|S�2nצ�%���cql�غ��3��`�C#3��c�##�����DA�v �T��0��m����hCB,�ja��0*Dba��P)*ވ��6D�J��3��łE,�(�k�Q��M*Uh�b��(xm1Q�xL4��8)�-�q=�D�U^	�Z�$��hX�c79t��=Fl7����|"Q�JFa2i�ȉ��b:���Xi�t�T��,T�:���Z��ֺ�lCx�����^�ڷW������WL�K��R׷�����~�;�	��ED��{���klZ�N�6ޕ��|�Wn��҄`���?ab<�1����?�hW�ҦbھMu>�*!�T���o����~���;�ۧ@�����3,���>��0�:�x۰�r\7�NV'�Z�? �͠���
����_Ɩ4q�B���U��� �2���d��d4���%�ii��K�6̎���b{k�j8 ����V��ʌ�l�(�#6-!$?���p� kS��������ɴY#8gp��XF)�W����s��G̎8:�&�Zr�zM��ve�>�a�g���ON���>���?�<������Z�=�qw�C�F#��qVY�,x�`��~��s<��|��lmn ��m�x��2�s��}��?����G?��G0��(����cBL&��P_Ӵ5w>�,����W���^bs��h�W�C����#�{Ɠ	M��=>��V�������;n�y@�JWR���ʲ]�`���ɐg��A5|��xBi�Q�BY���W���z��\T�9ӣ#�}�O�ٛʭ[�0ư1w���	�13��9��#(�儹�������G�����l�Lp�b5⌤JJQS�@��h@�*<���(���h�����bkk���.5bE�h2���(�����-�_�H�ث҆�mf�/�Rc��f�����Q5����8�1�oC4Xi%X+�x6��v�q�k[� ��5
�p���'�W#XREK���FBT�i	�k�cpEAT]�1�h�����)�����1���1��dzL>[ɲ(
����MB�iN��(���H�(�����<���x@�%eʧ�4���S���7��z~,�%��9,�n��e|�ò�:a�h��l*-L�Q�vP���I�K��Z�����z�1�V�ê�6�Ν;<��4��W��\�uӨ���=����,��* P���	8	��X
��Т�Q/g �*b�6��T轡��?}�M���ݹĥK0����/�ı>������Y���9�Ұd�q������3}����`��Ƣb��l��8S�6��W�����p��.�I�d8��-A-�i���m�߽�dk��y����y�L��I�;5)�k
Ga,�+hb���X��eQ`]*AU�m��&c2�1� gk����7��$���>g��{o�YYUY�7�E��Q�Ƃ4��@���������E�e =Λa@�0�a��戶�#Q$5����ޫ�����.����q�fV5�ZlJM�Hd޼Kč8���~߅v>���y��[���}R�H���Cj����Ϻ]���ϧ�>k�����c���p�Z�72�u$�X�����֏���c���Wv'$o��C�p��G����-��7����+Wv0�,}��R�m�K�����-G���4-J�O�_�am�)ʂ#]��t��PJ���q/�b	>���������>MQ�� �cL�-����}f�1�g��S�y|� �uG���Jcl��N�|t�.���w���b�]��R�Ӑ��R��/'��X~ު%�Oz�R��,P��5����L���>|�xTR%ZChm�$���,)^|�y��^�g���}k5"
���c��'''j6�G�Ь���!xΦg�m��S4vL�>4"1�I"��Y�8��ql��P���F��Ry�4)��Z&�Y�I	b�q�齂5Z[�Ŝ!�k����b)e8���^�1I��L��
�"Ď�d�QS��&��cDooF���~�1�R����-_C��J��q山*c����,ӧ,)�?/R�$	��N֪�bAb1O����w������|>�(���q��5��L$v�m=�RZ��{��ۇ{׮�ͺ���Փ���*����S��[���~���KӅ�c쒮�Wj�B��4&��Rk����#�e'�%�sw���$�a�i���}���4H�n������h������2[�ns�ib5���>&�|9�S*[�el���i2mC��I�����dl�}��aP�p�7��˽ֱc��_�_~���]�a�V2�J���ڶ5,�sl�c&��{�y~��W����l�R�y���~}pW��5Xm�YJW%�B�ǐ�g��aB���8g|$dQ�����kLF���~�Ǆ�e\!� �V���$���Q�iړ�u_�>��.�o�U�Fಜ�z٠�ؔT�АT��<Ea��-'�;4��t�l����?z��+���r��{��o�?�/�e\e��{��)�fOX!�.�ܑ����]�����]��\�5�_�썶�F%���:3}C���pŘ���[o�g����{� �|�J��y�Z����)�t�����%��]gsm�����h����,jR
4������~��?���Kl�<v�O;.ϯ���mۢ�����rQ�K��sy|�s���{>{��A_�R��g,�9��o��W^��g�ak}�_|���66��>���C����͙˔.��E$,�?�E�0;;e��7S0�L@ �@m۲����%Qʠ�,��Ƹ�{6nY�L) 1� ���t�A��kT0�0T줘mHR�������A�)k@�����rp��2lF;��,�gȃ
B�������(M�l$�\*5��5]�0$��2dKt��yã�]�o�s�=W,�;�FS6O�èIHʙꔲ:I>~ou�7�DT)�W�@"=!�tm��	Nk�LֈX�"��+���>��i$v��cR�h�"�d��y�~
PΟ���Z�f:�L���l�b$�K�D�T2�U�2�s���灐�b3�q�Z���l=�=��ؕEŃy�G��r���X߀Ã'3�(��U�����=8s|Ri�ݡ4�*+�XIL�@m�ȡΟRPy^jX����Ӷ�c�D�(M�\:��a݈�_�%����x��g)�����SG���7�r��u�z����{x��S\f�����Z)S8�����=
ED�mA"���\��~�|�����o�)0v���-^y���%�D�,z�]��	�$$��3l[[[@&E5M��p\�,��� ?����������MI`�j�DD��"���[�u�l������c~�_�����IL*�IM�g\�o�X���e,�AE!rvẋ�}��]q��1ׯ�0����U���m9;;�YM����;��֛|��m���ZML9�D�
�I�tDbJ�2�[�ܻ��ݫ�nl�QtmK0��D
M�/<z�����cP���5-���m�t���@oU�XfE2p`K�ד2}����c�����o8ހwW2em��ս�vm�/�U~���ʋ/=��x�o�I1��r��=�ܻ�b�@k(]%9��B�U��$m�b���6@@���uH�h�~�$�L`L�<��>�ڈ&�{v.E�ҽ��ܨ%��h��!F ��V3�0;�^�NK�z�(aI�QY�{Ũ@kM��sMU�Y��UI�JΦ� *�K;���ͥWb��A`J�y��HKJ$���%��m���zi.��/�����BΚ&�
D�Z��lS�\�>Hv-�]��9��$�m(J�-T0�E��Vִ֕�n��!Z{"U�M?x����x��:��e�ү����Ԡ��͛�����b�C	�AL\H�_��!�����hKf��eP103�Tbvn�j��c:�Ҷ-���d?ĵ���O����k~�7�ĵkW���:�0 �(���%�U��<Y�>ڶ�m�eve�֨4���	�O��}R�OD~^��}f���$��߱�q%/��2�<�[tM�qt�iy��*�:�X���:89��)1�H�cz���`M")A�6e&�]T���c�ꀖ<Y�$�63s��1vFU��`L�}T�5���(]v$899�n*���&�?�V�K��GW]e>�������-��Kr�R;2�~����w�XD����K��`lD�fѴܾ9;����Ӈ<��#���8;��RYJD;K�36�Y����	�*)\)pvz̷��/X[[cT� ��>�)M�55)vLώ89="����x7�=�_�P�Đ��$�ȁT�8�rx|���w(]�����W ��wl���,s���>����$8mxZ�Հo��2(*(����kVE�/��e��tP���X
+E���&�W���˯���̋/����6�-9;;���qp����I���5&eE�,��@d<Z��J�F2.�g�Z��k�L�3�z��#J��l��[�M	�Ǣ��2c�Gi��*^)d̲��#,�g�L>OԋŅ@{(���R"�\�,sŒ�R�ݘ^�h��J�Ϥ���y��R��#�@�ۜY����;��R��,9�Н�\�09x�1,�K��u&� ����H�
LH=�C+��ω,-�͘��H�A���%���)�K�9��DY:�Q�Zg��h*v��	=
^TJ����>|xT��u�vۊF���*�u�֧}}g�!��إ&�i܅�3]�"�EU��}��2�މv9Xr����g���2u]g*�����Ψ�*�y����`cc����S���vy�X�s|R�d�<,�]�-%^Vu�T�da�ՠo��w�?ia�y(�B�陼�īuΪ�!E���v-ڕ����i��,������ѣ.�r�
]�]ؠ�uM�4� <�b��{������*V	��k9����*7�^ac\H4!g1|��NV��*"@� ����~�V�����������}�ٽ/b[�Vk�*9���В��[X<M�,    IDATsF��8�8:9������\����t���+	���f(m�L&�D���Vk�V9!�-��&�LP=�H��ZZ�*JRt��Ih#8F;B�X#9Ќ�A:0d z�$��>�(�)�����k[LPH�>h�{�M�u]c�f\U,���tX������2�N�J�����q��K�����R�i�6��s٦����g�ʾ\��\�C�h4b�^x��ۿ����Z>��>��0����՚�|���!ggg��_�%B�fQ�PJQ�%�;�=�2�s���>�	fYB�{�lV�]&]��(3��țݔ�L6��~c��>�U<k�D2FDHBO��k���s�/%���(T�	1�e����k=D����
�!�#��uuX��\-��1��91$߷�D|.�O���,��]:�Pʀ���S����fx�����x<^�������8 O0���!�{҇��@� an�B�����6ڇq]�ηm1_̪���ַ�_�㣟_�*��~�c��F�I��!�����cӎ��*A�.�S�똢B�`�M$��Bk�B���g��ʸ������.N�q��w1�G��2�89��sݱ������w��z��2��W��g&�	Mӡ�FG��:/�� 채�>�*�y���I���}Q,x�)�H�<�&�e1Bk�'�>0��:|�ΒR�M� ,�g�pq=�M�1�@Ȼ.���b�DT>y���Jڮ��c�J��H��q�1d��s�%�y����/�)���Oh�\�$?�{*�	���3l�bʒ�K4~����OL۠;ێzq��?x�޿���X�1�ٌ�b���,�3��poL� $O)�Γ�q}prF�����f�`R�"����R���0�Цb����^y�����^f<���#f������c�+0�X�P��Ԣ�`��k�$����-	�Ǩ�C�$�ypvL�E�WH��)���s4O�߫Y�լ����l (�X5��Hm�H�s��P:au���)��d ���\���Y��:��u���ɪ y@e����'_�Oi.�����Y@2��.n�FG+/���� ��~�dܿ0�TU@K��[�������5B?R�c�B�R ��M����W�,����{����Q��>���������Q_:,������Xl��q���{��f��L<�nnKt�IEI���Ǚ+-h)ʼ�w]ۗ\=�����lpzz�3�).���L�6���ec�2C>l�677���㥗^�W^a�ǜ||����CX���98Q�tI��ͥJSN0�-�1��Z�����欪*Du����r#�Y.����pơ�b��
EL�D�wC�pe�[��)&u�q��K��&0CP��h��%��r��N[�3'!O�S��F*��O����=ñ�y����uJ	����r$��$GW?ؤI�8�|��1�D���i��}�����ID�d{�e���$��j�\yC@ň��|�R҅V�`��U�k3�ו�pvz�N��֞NO��3ƚ�Y�g�y��=�'-�Jb�����Q�S}7o�L7o�q�ԋ��AI=�L�!	>D)G���$�8;��오 %�C�	H�����䄔�E͇wnspp�h4��8<:�J)��)u[c�S�~�m�����3�<�̦���1��!S��]x�J���jľ�.�a��ߗ變���!ڶe��.'�Ld�����i��6����Bz�=vy�_���b_��[�@�<��rP�:��@��.ι~�]>�{�G|������g>] �6��4�C%A;Ka,I11oj�6(k�AR�@��i&��gM���&v�7���T��d�aM�i��zA�,�E��(2�ue������Zj��&���������o���D�2c�$��z����R�$�p��h�$��gQQ��(ML�#���XC1Ҙh3x\G��^J!KH��AZd�hⱅaTd1���������)un�vy~��۶���ev�m����M���Ӵ�VU���ll��t:�����9��������UU1���2�N���9�������9���@Y�,[N���H/�;��$�C+�1M�\�T�5���!B*M�µQ*c�SPK��2�ѯm������,^9Ɠ�<{Ѵ` Y�b I��H���W��(�Z-�'�$b8ߘj�2�^�4EAY��ev�ϡ�+X�,�f��H�xR���������D�QHt�H�.�XIT�c��pI"�:�$&�5�P.��M������"�����J�$ҹ��l{29�R�#J�[��O�yL]gT��k/�S����w��(�V|S��1�&��t�]B��ipe)1&e�5�+2�8�Z�v���$@
W *���I֧�֖ʍ�WUf���(��o�������}�Y������1fyc����KA�%-�U��0ПTz~��-�N���?��؞Y�rY.w�s��A�H.�̯�S��L������3��"�i��\��dw�����9>�������T� a������os|4�t�;�����A�+U�Y�͢fT�\3�k2+�B��tG�����A��L�ߚ� )0��Ѩd2{Weצ}���C�/K�1��.w��)�jV��ṡ=}�XeI�u9�c�J�.�B�&I��8kp���U~l,�p�a��jC<�u�"^Z�}X�v>g���j��	j��E�l���A,ZU1��Ç�<�LC��UÆ��nX�{X�>�~���i�~��KU�O
���Cw</m /�_��|��5�ס|<ظu]���׷7��Tw�&W����&M�pxr�$R����3��E��mhЩn�&H@�E�yO*�ULA^�R8OzĔ(�k��Q)bL(ՓP�!��+Eˊ�P����}�ߺ��A�֚�u9�3�a��ƈR�IU]���ka^g����>j֞a��r=��X[,��(���\��g��\�UP���(P:o���m�d$%�E`:�+�-F㔱>�wI"��PS��Ux���N��Y�1Z�L�ԑ��Q�BJ���4����8c�c���AQUGhӖV����%^�w�o׋B��>�%��hL|ԺU��wQ��s������w�?zp��Ͽʯ��o1�w�fZ�I%Q"����.0.
�Γ��gKfuM)��x�h4BiǼi�ǜ�f��_���)W�^�C�tX�2�vri������3}���Cv�I��1���l��/(�vZ�#(�9��~�kb̯�:I��)u]/�1�=���ǘf�%����K�x��jИ��^��������&��[���g-��Z���K�so��]We�����9��BYE�	c���	�g� �b�T����U�� ���F��>upp�|:є�q��с�DY[ۦ���Jn�f۽m���U��O�\���KV�gi&���� ��v66؜\gws����̆���}Y�˟aR_��2*�Dl��i�(�
�
RR�ń���L�
5Ei�!��g�[�vX]������{�?⭷�����dz{�4d��11��$,�?��w���\�/��Ļ�T�6�K՜���0����d�����bY^�_��<�y�2��:㇇
� ���0�/�����z��l�9����|~ڟgp�4I:�Wh�PJch��}3� _�����:��F�eY�)8�L笣g�d��2�A�F����g��� )S$a��$�r�f�-�%8Pl��QYĺig�^҅�PBt��b����F��8|����eц�ۈh��s	9j��eU5��<r�RI�F"��)��ژ�� $k�Kb�(ZDy�@C��AsY��A:��� !�4e�C�uRZ5��F?&Q *����t�Gڮ��,�WZO��b�>��?9>Y�����uk2�|tvv�nݺ��������o|#Z�tA�mT��:ejچv��Ç|�{�t��ʫ_E����5zM¡mB�'��l~F�8g�eMΜ ���{��Xf���&J)n߾͇~����:��e�(1�zͥ 	gt�>擤/��S����o���v�)KCJ��K�=�G�L�ǘ�a�{"�Tp�s�]�y�
/��I��j[�S��˙B�;��h���N���1>Y���T����J	Lv�2���+3OR�j�h4b>]d����&�H[wh���V�R��O��:66��~�W�\��m�J�A�Z�lIQ�K��#?��yd�(����]�|:#t�|�����*D�Y ��(�}>�W�y�2T�o���W��	:o������.���U~��x��u�no���Q�rR_��iU�a�,��/7��F(m���^�'�6�����A��e�ch���܋/PM*O�xx�0c1����z�]�k�r��t��_���փ�k�Xt��@�B�y����[Y��*���`p�?�[x��o����:�Z��1�u��Ou��lvJ�4KG��k������nBX�Ƙ�n��huf5��:�?SBʏ��X�eV|r�tV/��j�`�!f۽\I�Rk"BL:����%9��1\3Q8+h��&��ߡ$W(4]3mU	Y1YD+���0�(�E��*�yH!%���䌨:�&���耊1�d�$��1��Je�B�Ť6�W���c�7�R�Q�R?�H��� ")v1�n4��z�4I$ň�DItZ���Q�F���gWRRJ�N9R�)�@�:��EQ�RJ�`��6`���F1���c!Y���=|l�����R,�v][We�������#�M��������NO�)���͛	mۦ(ʏM<⵱�j���x||h�|�Mv��g����]��DaQ�����ʢ�����|��tF�����(f����e�w�L�X,|����w�_���q!K�m��檧��Rͽ��0{x4-���'v=��cT?��ˌ������w�mH�L���������K\��1/�D��'�<�W�.�Q.g
����Z^�y{��Y��N_q���1�Q=z���&k#�ɓmU�h����d'�p�j4bwg���M���I1b�e{k�kׯsew7{��`|��{i�~F���ǿ�5=z�3�6�еs�����C�y�������>�ڞߣ%�xe�	)���|�?��b� ���3}	MJ�-*����+_�*���*���6��u7$\,���q��φ�M1�2�"�{HP7�B�P~��ӏ���@��w�;Ϛ���=�}�y��w���RYn�e�>��>�|?G0��U��g��n.��9��Ԭ�hV�g�˺��dyNC�ou޽,[�j��Im�����ܝ5/݅���������_���)C}:NNN�������l�����X�0Z���Y���|���6%"!%��m��`��$%ڈ��5L2F%AG笏	�V��*{�)QP-� ���Et�f�����[��$*DD�GR��9E�,E�����:�R-�)Af�譈?NAG�t��L
!:e;�z�/Ԧ��h�{�:01F�I@2�e�Jr��Z�C,�1��ڤ�s1�co�E
��>����AW�R�q�I:oA�l�K2��Ҵ�b1��8U��Fb�֒��|�:b8DB�	�ċ�6�I*��T$�BE��`SLN}*��[��	":F��Rڥ�x\� �t��!��HL2���M�
��Sw�y������w��6��|��.����.�m��|h�G&���j��*�M��|t�6��o�M�s/|���7pE��]h�� ��X���1�o���Gw	ƕ�MM�;�r��ƣ��w��?������׹u�V�yBJ�΢�.�!�C���K$g&��T��x��d��^\�.���Up�jau��9�d0�l.w�������W'�U��LG���]�Ւ>N�>wFY�N�>S���/�X���rPk2Á�#m]s���x�}�]�P=�E�ޕ�dbFR0*J6��xv��n쳳�E<"���2��I/oQ��^��!@%�U\�v���u
��8���7x����[ob]����V���=���f4������c��Q�K�~��xOkB���#�׷��ڥ(3S�	-�"����Ĥ�*���9�yՒqh�Pt�'&ͨ1M��UD��ʡ�%r����MP��Y��)K����mP��t$��-�t�� �3<����'a�T�!����WH�l�;��Zz����������w��t�z�u�����r�
���<��KH�q�����ѣGܿ���q�-���$�]�-�"aHQ0�����^}6h!6�	��]�6�4���?-���v�)tSRH�ke��Ց4Ac�$ʞ�������"�nH�KI�Z�H����`;���`;��N����L�T�E<�v�B�Z��C����͛7;��7o����������YF3�R�r�L�Ke��t�m�Z���}-B�)�I��6Q�eT2R*�]J�������_��$c��H4��N��N�C��%%��(����T���1XM, M2�A)���D�26D	$/1��$m�^Bx��,=�����VX�'�R�(U)cJ��	�^D��C�����(�]�`'6�-@��zܾ��k�֭[�d2�����3}G����6v�S��o$ԕ�	�4m[�빤������������7��ۿ�;���L��P"XWr��>���ͭ[���{[R6���zu����$�s|�]�r���-r�>��7}��;�Y�~�����|C�u�f3���@�x�JXH��f��]N(�I��30}VŘ��1����񒲿X,��j��
�]=��.����0�(Q�}1�r��c�Zf����s�RFH(��җ0�����6�@�iY�0��[��g��W��E��#���l�<VVWJ-˙Z.�U����^�!0�1�
$v�l��W�L5��|����>�U�{'���ccc���X�M�_.�>1���-3n}C���w��7�蒔�.%*m)ʒ��9M�,eo��ˀ�+�,)1�ϗ:��"c�����ym�����F�|^x>f6�q:=#�fm}���/pew��x��rL�\JʘMG�.�*c�zŇ���/���6Ta�F�
�x���Pn,ن�v �V\>k%d��֋Ռ_J��O�I/��h���s���>�^�h�y�l~��"�*
Wa�Ba(&%����`}�J}�O���ƍ�!&�x��G��sաq������x�"g)t-:"�4��3��d�>�L i�L
t
AGҺ�`Bd+A����I	�(I��1�h|��jQ>h���n��u1.?H]���k�(#���o�{���{?=��o�M;��IXخ1�ģ��Ye۶momS��OZ�N�k����h�8��W�0A�^��A���(���l�>�N���D�2�����$��BҺ��!im,ؔ�7J�����	ګ:�dt��+���""��:"��d�j�H�jD�����dc=��1�%�-7���a����0����<�G��>����۶���h#���;j6�����GGGR������|����g�͛7���3}��ݓ��BPb��]l�J����b���,f���G�l~Ʒ����s�/��2/��_��Wi������_~������t�h��u%m�b$��'�����#&�k4u�n?��_������]<x���d�`:�����l6G�Q5���O��Z>0=U<��[,�e�b�^<	�
�&bub(˒�|����d�s���A�o8�����R�X��놅�9G�$٢��	i����%��i�[c�f�R�=(��m�msV�y�-��tߧ�WK�O��i��ӊ�|�5��|�<�sד�k�
��8g�b�ʒ���Zm��l�0�,�:fӆ{\�,���(HQ�7-՚�Yٽ~b�(
�
�vL��''��*~����u&�1g�9��#�lsT7�u5���=��v�$�,	m̦�*�G�N���V��C����e;D��"!$f���`s{��G��;x�w�}���m�4UU�������b����a!lb��Y�k�5���3{:y��9=;�l6���
�_���wx��W����_Ѕ����[lo��}�m<�zE�hpnDJR@T��������S����.�~��=F����2v�r��c�\��kw�A�]n��q�u�1��ʰQY,�ι�Fί��z�j����������3�O(�x����׾�˯�o�q�۷?���^0����sm��    IDAT��Õ5�*{�lf������Y���U���xD�^�a4YG%�(�����t*v�(U8�.�+��קg���zWD�[ԋ��h�����uR��E�I	-J�I��:�3��%CM��E"mЁS�T��̕R��:��i�ME����	�ES�H�֝E[�u�Q:c��C�����d�>�w��ƍ��t ���tW�Wڣ��SE�(ڮR�.��Sl�N��F�I��騬�$�7:��ѕe�&���]���@Yy��EQ(����Z�ԳL&�|�?����1��R:�=R���c[��h�(^=�1e[����.�2�m�˿.���՗�y-�z���y�f��?��{��{I)�I��^�"���o��7oݼyS_�~]'�nݒ��뢔:�_�D��g
�nܸ!'''҅YD���6F-�Hl}}ipP�Řӳc~��-=zȽ�w��	���r<��v	�C����� ������g8UKf`�u��o�{�23��/C��U����Ռӻ�1 ᓹ0����m�Ռ�j���`�z;�2�0��`��kX����g���y��rPt�=��)�l�_f�rИ����8������m-:���rlݓXW�9��FL&Fe�f�_�LҮR�eT���Ễ�Z����Y�(���p#p���!��5�D�Q^~�+���qmo'��R��jD�\^�,����Υ���*����瓼J}ILe�Ӱ�J�
�\A�f3�Óc�z�-�����0�N�ЃA����,��Z�2�K�
?ϙS�h���"u3�mj�7�4�C�tݜ�4G'3NN�\����~YS����[;lnoѶ_�%���i2�{P��E��T&(��ڹ�PyY-��*\�/�jyx��q��Bsf�Y�c�7�{{{���s��RJ����0���e��5�}�Y67�������N3=�sp���GG�����M�)���r��m:�2��u�s)�(�N�ֺA̩��$/]D�7m7&�p>��a�����]���C�d:%�XGm�B֊�l������(������H��;���1&km�˔�6fjִf2��Η� �@g��Y�gG7n�P����������ɭ�o��o~]�c��y-���O����h����qP����p�{o�븷�'��$����w��ٸ���' �׮��\����]������g��6����n"J)�7�P���������͛7?���)�X,���RlD'%)���(���$�o�D��}ĝ���޻o�������8�k��Qe�ۚE�bBi���v.?Q&g���
���{w�����RD[CL1냹jI�0.{��<!�A��qy�_� ��eЗ�;�hm�'�:R�e9�^�����~�iJ	���P����.g!WI*���I�ße[e���U �OlI=����+�(H0��'y���Y/��'��y���]}���V_Z�,�٢��8WR�2k�T�ƣ5l��7��D1�1QY��l]�!�^�[����9>��Y	���H)��_��:��rA�S�.����1]����J���~�o��ݻ?�������V�uF�k�;�`�B�\��|����<�Α��iO1�a�1(�����^f:��d��o0�����C9�I�h���E��mO�k��0�\� �ɛ)�Կ,�b��[�E]%nmu��Z�}��.��������[UU���q��5ڶ�?�w>� c�Q�+ƌ�&��g�n��3���w�srv���U���_���g���Z2���G���T�k��{�#��]�1��^z1��W>%E���
>mt!mn͛��jT�%��֣���6<x�+��N�y��jp�IT�Ϸ�op��?�� �������F׫�t}U�8;;���}�5d�>Y �)��g?�����7�xC2�J$��Q֤�bL�ֽ�M���1*K�QI�����p����[뛘�Q�����9;�*�0��l��*�NO	OY�Q�}̥7��!P���|��P�a���<z4������� J�����뙩)Y�W�=&*e�-ԋ����A�!?o��-�x�ؗ���x�s!C�	�P${2�~`�e�J�(҅�����h���^ �|�sQJaz�R*gy���������-Ύ�LOg�U_��nllQU!>��$^�#���\��*C&���4+��
1�",�b<-�i���RZ`:mx��i[��<IV�|���2�'rn��9��z�ؕ�>E
��(ʲ�p���<zt�ՀQ��DSX��sy��(����O�*RRH(�}�3P�&��FkGaRL�$c�E:i�@Y8��z�O�l.K��-�ۜ��E�{����AJ��b���1[��e\Ul�:�O�sl�@��d}ס5M�o|,���lll���ѣG|����3d:������!�����uR�|�+����a1Ei���C����޻��7�}���3f�:ox1�6�c�(KYU��UaݾR$��6!��� q3i�̨��iqf�']�����a��n�͛���-�߻�JYU� ���w����g��q|LpN��"u&�h�
� �����h*�-ZB0β��F�����@�+�J��q.��*�J)NN�X+6pz��-�T'''(�;v�#m�E���O����2鳢Ö%zE��w���%� ���)��y����TB���%&��5A]��w��%>�]��]~n�g�L&�e�R��%i���l/L`O._|���P���"*�%Ԝ��F�<HްVe�h4¹\�H�H�@MR`KK5���� 
��r�o��\�g<8;ʾ�"�q���5�5-Bbzr�b!�Mã���[o����%������tn쾴��S.g�SʎO"�|^m��}��^�AeW�k|hP��h�$!� ��e�TE���d}}�Q�G<XMu]G#]�)��͜z��ʻ�esͱh:��
0��Jh�Qo]��nyl�5�:��>����E�{�d��?����8;;���l�m09����{�fY��L�Y.3�m{,<")I�I���g�{f�4?�����1׼��ŌbbB���H-��I��-�f��X�UY�l�� "���Q��ff-��{�w�I]׉&�U����7y]����#�ׯ�tp�.���>�p����c}��tzH��3�N\�e���C�ܹ����{�pzzLU5vGتi��`�A�H���hă�cbJ�G�x^!�Q��NC��EuX����Q���?�<
�|j@��NB�a}t���ѻ}����|�HS�	O�ƤU<1ZF3�/Q�����R���x<N�u�\I ;m��9��Ϭ�两�\������,����O���R�g�.Fp�c)�/ט>����jR)�(O�վ�h����%ދ%g�� �]خt���:o]�i�T&�d�£���v�.����'�ː����^`�Y�]Ӭ��Nd�MSqr�`Mz:f���;�(
��1{{{���S�z�xx\S5�`��+��ٙ�a��,K�����O��_��=�Ō�}���)���%BF��P��o�nS���$t�o�\)E����8�`]IU� F��A,Fl�vM����ʵ��'�le2�"g4����d42�QB���89z���}�R�p:]a�!4���\K����I�_�1���2�ߺX��?�?��:�,ĨX.�<x��g�]gT\[$w��2�֮!0�5��)[.���ײ�i�֐��4~-�������,������l���	�gS�k�Z(��kCʸ��2]�MK��v5&�8�PRJ��PR*/|�Jeh\���'d9�9͏�<���N���!�\2��9+���-uJ�k�����yCp.�]��191��X�d�\�Z;�L��%��9�Ʉ�d�JFy� ��j��I�n�8��5z��)K���6 ��������^b\��&��D�&Zǣ��me�mj��-�|li�2�I������j�|�Iܔ�~�Y����}��q&#D�!��uBЈ)˒���Ez�
()	�1_M1�0�p��^�����:�@�gU/899����_���H����P�9�k�9Ҍ�ӓc�}�!}�!W���h"����2��dNc�o���~��~E�����g.�\��nb��`��x_�l��p6)�Ȩ�J�ɜ����	�W�GH�qu��!j�`<Bg�|o��d���=2c��s�w�p���rNc+�/h�ckAA1!�;�kZ
�wTU���@���[�D�x��:~� <���a'y���$��Ln֊���u�8:�������J�RJV����L�S�s\�zm������'(m8=�rt|B�8�T\��E�L�g��2�� �Hcc�Z��I�=�Y�j���*�R"e!6RHʀ+�@�΅:��%��zj�Ş��;::{{{ ���T	�*��2� B�	`�~�i�7�c8̑��r5c6=C�W�itk-�'5
�R�}U6���a����畗^�,K�?}p{-q��i�t�۬�I�M�ԙ�ni�;s/:}��]��8����1]V��j�M:�"2*NϷ������$��R
緛5:G����OB�O�������N�O�=���c ����ϑD�b>�SU�)��i�b���LF���|�;o��oP�%���ܽ{����/eN�S����#v&;g�������G(�2����lN�in\����1�q�n������'6�9�_:���L�����8�D�J� �)ڌ�a���8� Z(23`r�͛7�Z3�B0�s�sh�s�{��x��!�������x0����hA�I�$!Hf=߈��Ĺ��ŝ��S��~�ƹN~l#���]]� a~7JJ}�Skm
$~��}~]���hKʉb00�毢(BqrrB�0f�d�f�u#���!�̉A`��65B2��,M���R���qȤ���h!�*�#evp�ɫ�<���yjP��ʻeB;'c��e,Px6Da��%�w�P��L�}�&ZJ�U�'�%:�R�I<���Q�3�_2���]�>�`4住�嬪�=|-��6)cb]D�ClB�'��rI=O�����
���T����đ����k�pEA��5�sG��F�v$��ш���ш�j{>�Q��Ӻ�h�}� T��ު�X*�x����g,�(4Ҥc�
z]�k���ڲ��l��?�l�IEuQ!Q�(-p? 8�My8;c�sA=A@f4�ȢT�N����⫯����{&�n�w��#n���g:;ag8�����OFL�ƃ\K�.�$�!2���|z��l���c�,c|x�Ji�޹˭[���ڿƠ	T�$zEt��j�z����mÑ��T����!��L�a!*�9D��	/(�%�@
lA\�`�O,��rF��x�9?�1�FL&4�������r� %���&3C���hF<c�L‸X1/�I���,�r�w�s>K�hw���H2r)p�$���# �V��H,�� �D�$b@����}ָ�3�!S��@��Q;Bw��5���0���|�n{�!���$�bIPK�h�*�W�*g�<#�y1g:}H�^چ|�SN�����BtT���e�(��b�S[O�
e
�R�& �%�Q!��3Bt�:˩}���=_��tӃ�(���dY����D$���HU6��n�7&j!ڦ��$8�ɵ�6KBY1���<�ލ��[����-�Yt6 �o��&�I����q�h������ ���"�k����f3vw��9��)�$(R@���]`��3�ZQ�"8�$Ǧ�J�DV�Sޛ�L&��^F�U������ů�����6j<��퉝>S��j�@	UAH��&��QV8��*z�7 �l�	y!"o��C���minUUF#ƣ=�v��ptt��cM/��nӤj���\&� �H��������~��G����˲�����k;��.��W1������$v�4������Ͼ����7r|�z!������CU�h�g��Wi�o����ۿ`>�!�g0�����,�GX.��eI�u����h{��t<��5�����y���W�\9`�J?�֯�K�])������֦_L�9Q��4�"]M��ԡahr�a��8W�G�4�lg�f��{���U�9���W%���e�bV/@�)vwǘ�yd�ne��@������< ��Z��)��5���p.zdLk�T�kc�U��/�kO�5y.@i��8"F$�t�<�2jv�;�U��p���b"�il�ZЙA��R�Ň���<O��>&̥1
$R�q"uR��ֳjV4!$�J-1m�'Ĉ�ms\�ԫ�S�YZ/BXBk�R���;�p1��λ���y�|�XϷ���l'�"��2\�e�/V}��ٛ�s�9��9���l��Fu{G����kmn)H�TQI�P4v���{��2��T*SR���u=�|�X��ƞ��{���ѻ�
#Dp��"�=+df�RB����E1�v��G�m�VӀ�bU���!5e�%�.K6�N9=�1�9`<9��uP�����-�K��[N?h1֦ITV˶SJ�G�G'R���1�;�q�Y�&h"���7h�Q���d��o�
ߑ(7M���ҿ~����E�b+wU��e �/��ߙ�����r	@����C��������c��1�6Y��9?}@9��*��\[/��s��"u�M����s�!0���4qgH 2�s�R͖�'D���;�sX?����孺��;��!���!�#���_� U@�
�'R��Uę��<n$�c�ݣ#~��[��V�ـ��T�"g.T��̝qڜ����n����oeZK"�y��-HŰ0H�	Uē:���⃇�2�)��C�����*b���$%�%F*D`A8I��Z�:^U!p���T��(0*���A��o-R�����c�Xy�SW{�]&�<��B"L�.Fh��<;OA/��L4(�Ur�$'ELNgHN>���1�!��svww���[+]����0�۶%�W��3���4'�1���>��#�=���N�&q^J�W�\a>�o�/Z�p�{�/�n���: ��ɘ�k!�1D���պ�
̞`�>�/�=Y���M���>�D�;D����2u�n�)SYJ�&L7n����:�"DWR������J.g�3�=<b��u����Өk׸����f���n�2��D*R���.�B\�~m�bv�q�C"�l�1�7�C��2Y�l��Ď3*�G:GNF�e��+�/2���:c}��kj1Fc� F���>��s��l�[)�@lȆH]-)�!�������=�����L�����{Ì�ܠ��0��鮵�婔!"�\s�3"��ݻ�99:�D�o<��ݖ�$�V]�b�h��k��󰋍6�c�����XD�P9�,�RhS�3�E�+3z�`0�Xc��ݵ|��?e�w�����7<<=&�$��S�{9���fF�*qN2f�������4n;\�w�,Ө,G��sM���yQ���GȈ1)�Y�{�Uĕ�L*���E�"ϱNPVZ�LF�lE]O1�K�RI�\L�EA`����
�R8�q.2�r������n�geK\��ZVh�8�z����gܼz����h�T�� ��#�B��1zD���3�߿���C�޽�r�Ļ�]����k���w�L�h�c4�`�?���>����E"��ߵ��گ�\����;���;==�z���A����
��ړ:��F���� |BHC@��b�O9|�ڗԞ��;�ʙp��Ѝ��P"8?�2�w>F�4V�V˖\�я�pg��S�?@*[ "!RElH���p�������egw��xD8:��kB' :�#�Τ���z���э�bf�_n��>�OLj�2e:޸@rchg^��2��B7�;������4Z��t^��\!e���n��2��{�H��Oc����6*+��	�Z�-8���9<<\ӽ�"�h!�D"AK�̥E�ͺ���+MUr�{����!?�J���{RiI��*k����R��������(�!�UJ!�GI�w���`2��4(��%"8p�ipq��5Ŏ 7�|�
_�����GGxp���3]���?����P�cM�H��=�    IDAT���n�xE�Tq�o���ɇ�̻�-�Œ�p̍Wy饗�FL&��4W�V�")Y����C~��=��KY@�^�C �A#<s�Y���H5���6����bIm�i͔R��L��2a���|��_z�o|�ufƭ�>��_���B�(W������[���;��<����
�Uհ�b�m]�3��Ղ���srr�·=����C����5��m!�5�2�w0���N�[�_�H��wN�Ex��&\�)�J��ck,nd>����I�N��.�~�����w|!v�����	t�&:tBB�T�A�����}j{bL��	�BB�2	SB�]#��!Ɣzvn��]��!�=e'�.Z��$�R�0��Y��g=<e��&�`��h̕+W�}�>ժ���,Z�.�D��k�U:�ۍ��e��Ob]���m�#l�`�d�Z����u����T�.�-��w�w?��]�:%�v������וտ��9��Z�X/��k�s�fZ����~5u�VU�b���Wc14H��_t���!il�Ķ�Je%dj`�W�~�:M���w�t:%��r�D�D��[R�.�'�6I��TyW���D@(�(�D��A�;��˯��3�p��!7���rq� W��8?=����4u��+�1�����������sL���e��Q���[�r�`�Y�)_���>�xƭ�������M�1�eXBT!q>�\U�u�x<��7�ÿz����⋘�%ϳ͜��� ����|�o�zĭwn��G�����`4d�J�@��������J/8:����ý{�x��!�yb[�PR&�h�B�и �������o�g��n�,���)�����#������_{�[��_A�@��� �4HA��פ��5:ӌT��9�{W0ِ��-Q
N>�ڲmj��`	�!Q\TU�^_�u�v�����ԕ�ښo}�oB�]��l=�W�9�R�u����-�-��sP�ր֤L�חL�U@MgS���2�H��1z���O1t�ڗ؞��[,�x�J�[�d�B���E7�ʄ��.�'b��%��s0���	���$i�Ve����墂��b4���g��}��%�ѐHj��Z���i#X�kZMδ�zo[I��2��i��Mꮬ�N������m�GR���jM �9|��u?myW���c���x���,��z���1�����S��;�Lf���z���1Bi�ƒy����P��%X�6��hLQ(!	�b���Eƈ��$(J��:�s�������k�ٌ��QK����r����߈����Fӧ��z�I�� ���_��^c�`���r5%�$":�w��SN�ψ.�O�|��-��w8<�x������7i���${�=�����0��x���woS�#E�ɖ�����<��g1e�����7���7��������?�:�u2"�@L�m!�i�L6��3Wy��7y��78ؿ��ܾ�6 *R6�*�����+<��WPz���Y��o�M���3�F��V
��6D!�A u�x�
Wo�ȵg_�@����F#��(oȲ���.��(r_���HzM����AʰY穛����:��/�3�"x�ώ�!bׄ���s�O��W�Xc��*��u��sY�o��]pĺ�#�D�}~w���n��7:���,�(����6@�؎A@(ك�D�w"����E�#j|X���a���G�S�C�'��9��P!(1�{�BJ����#{��׷6��ðvH:G��,"H�ሽ�k#\ erbh(˄1��6��nk�\v���LW��ȑ�#�-5u�nFD��EI��庝e���e�ēX�p�6jO���ڈsv��KY�����A8}�sk�{��*�n�O1�I�g8פF�Lᚤk}��+B ����x�͂I��A`2��/8�M�5�
��(�:�mf����HH:�&�_��8�5f6l��TЄvSsM$7��!���䭂�PJs��*�kN�Θ�N�Ww�yx�Ã�P�h����jQ��FF�_�kO#�EI��:{�Ƀ/��c��9�����������?��]��������8�B��H�(����X�\A��������A���w?��)v)kO�z8$O�"wv��wߢiQUMҝ���f�NNg
Q���� /2��9Z)�,#xP�h8�ȇX/�JB�$U.�w<�l1�G�lW ��mCŀA> x�=8�瞧\Έ��*�*P6�c���e�J%]�G��5���y�����.VQ��6�0m�O�܇�tkS��^�\(����1Ɣi������3�jB�!��R3��-R̤���<���?�?��O���+�R���e���4������j�r�RZ'-�NU�&�~��&V@ˎ=U�\���v�%A$��PIZ�5�����&+��; �8���2M��ʵN�G��n5{/k��;�}��s��Ɋ�H����}j"I�ä�a�j��!��/�[���b�.Cv1&N�~)�"�;�����6e\�"����Ν;��x��g���4���3�s���>�T.�]�wL����>���������>$)ѕN<B��nQ$�b������Ae)�!Yw�^�ʲ��:3�ImBH��&�� ��wB Ed^V�,'8:;�t6�iB$���b��p���$�k�Z��{O��Ɣ����-o}VB�;ɻ��I�`�eX<&����ٔ�����6��}Ϋ�(�d����>É9 3a�г{�%n޼��sh��46�E�x��`1���ѝ{���_��1]���`=VW�y��}�`�[/+��z~������-��9�7<����o�����v
$�dgr����)�,/�^0_�P&������cr��U�`r������hYq6]@��@�Vx-��N�.Ғ�w��y>����旿�%y������b�Kդl���.�:���k7��9�iq�����x�`�Z2��������֞w���_�;���]VuEVYFӤ�%�b<�p��Unܸ�����կ���Ͻ�p�qxe�����V3�R8�BT.dĻ�;��:5~�!]�֮)�֙�6��>im�@�{ t�C���u��.��e�������>Qs�9�:\��{C?�fah��HL�*�t,]0�g�iD�"6um
�����j�T0��� O��?{"��j]�s9Ep>z��QH��A����8��(�E�ڢh�l�ƝgKf�����}�$ӻL&�����,�+�!�QjHJ�z۪2�-�s�Zo��.ӷ���8]SDb��Қ̨��iA�En1b��`P�)q�rBQ�F��d���j�X�i_҆u��7�R&���p�^��uv/e(?^r��e}m���؏����?����M��M]˛n�� ���qHi���̴�w*�����[7�w#D�m`�/u�$���rU����w��9�fMC����v�I)%Zl�Mg���i��������CJI�$AIVJb��2���i�����F`C�ɑ\�Nvp%ӳ�Um��$b�sD�L����Ղ(���,�*GsAm��d�g��R����?{�-��ʟ��C����O�ۿ�[>8���4IUF	B��w�ի׹�ʳ���<{�r1D�{�7�{��^x��_���&F�C��@��!#�)��y�y�կs���64��,8��dʉ�(����'/,1��u(��)��[������W����LN������D;2�Ny���w��ZK����x�eȇ#�!"����g'�������q{m�,ؿ��}E����Y��,�J
��w]�����C$:����������b n�5�������i��-���C�R�*�-�K����#�'o�^�h*�(D\;-���!D���@�x9��B����_�1�D$�@���℻YN���s|������������x�x��;M]R�UXwe���EX�Iڟ��c]��=ן�J)��J
�4dENn2|41R55��$J H����qC�9}��uqx�����9��x�~�:�Ɉ,�Ę�SG�/m\� �>��!��E�>ٹwc��ߕ����9��f��
��0�nC�%�<C�5���q�u�y��y����"����J����j[�^g�c��GR�����Š���\F��T���L�04,WV����5���3�v���!r�`MRJ������Tu@G�S(C��b`~��;��z��.y� �5|>�˧����\�k��&�n<��|ͽ{�����G�߿�(˚�jh|R�@hL> ��q����u���%7���}��p���ܸ�?{� ���{���)�]�j��g^���9w���W���4h-[8�!D��Q&.��(��Ӗ?/�_^V����_��=|�6�|�@��B�3CD��<�V��lJD'꫱���L��A��~�<��V��.�-�'��n�e�,x��]t�.�/��J�����k������[��o�ɤDH%���k��я~�T��Ȟ�髚+"��EAĐ��ZA
�]Kbk�[��µD���'k!"	�sOF���h��s�j�o�x�����s��Y,KWS�U�4U"�\��&�`��,C)�`4m��M�[4�z�i�n$}�ņ�9l]3�(�K�LF#�Z,�d4�v�ȱ�>6M�&�����E�q���9����}�\��0� �+������r�.R�\�*u�_��u���c}'���k+w���%�&�� S��V���µgO\g
A���L��A���(|�px_�뚥�(�ϧ��۬�vA`g����}(A�w�g��甍�llt��Ѐ4�)(��;=!,O8��M�h�9���wyNe�H���+�-.�Qx�8Z�yx^��Ś,����p����C��`�f�l��L��QJ�1%	���J~����7��_3;?&�
�cq�������d~6���y����׾J�<����89:N�6F|��4D�� ���T�^|�?���y��w��f8QV�$�%E9-�xޖ��ylD�{D��Q��*lY��d4��j���$H�9R�hr��8�s�΂I�S��9������H��ҙ����i������]�8v��u�����u��e𕋙�K_�A�bh)�D� �U��Z
IPR
���R*ɤЯya��˿��ŏ��/7U�S���)2}AHQ�c�QDA�!D�Iʑkl���^k�u�.()pw�12E5K���)����W���=�����n�\`/EaA`L�p(�~�()l:e/frB�(�����s(18��&�w!A&�#%"�V��i��(@K��
-����[,TU�sn-�V׏�jO�uYî��{鵍��Ŏ��ǡ����vI�r����u��~8��l��A�ׄdj�%�Y�]I�����I�Q��J�nJ��9���!�+V��Ya�%מ���4͚���%�si@�yY?{��w��(|ʸD��5e�����^�
����3:[�%�����ūe
\+�pT�(}��5�l�K4�[�0�K�ǣ��h7�S&��^�M6��	��g��������;w�cw�">�4M���Q�&7�����;_Q���������q<����z#Ā

�2DTT�����,=�p��n0��?��?}����6�H#��k�TD�Jj1�ֱ􉛲�4��M]!�G�$/3F��B������f�'b�� IXJMҠ��B>���|k�ɞcwO�џ<Hl;�k-��!`]�K���8:�ʶ�ww��n�����\Ƙ�|b���wY�.����(��h�
�C����S��̞h�ԶNٽ�VQ pi�ƶ'���=w�9^��:\����������[bg)�"��>~x��x�`�q��3�	��ٛש��:[2�mCpĹM'U�	�w��~�i�JY�N��{]7QzD��:ӧ�a4`�%�e4��,	��(������lFh9�V�!F�њ�>���:���bЋ�z@�$�-��n�J�� ���i}��Q�sS����uI><Ew�!D��0��q5Fzr�6�P/��S��/"MU�Ɗ�1�>��V����od-^ꕧZ.��\�ju��ޢ��6�,�kb�����TW�o,%O�e���d����>68۰�M�e�29>"d�!�Т9<G�S��y�:�gXh�sc4�h7Y��������]>��`A��DR5�5��p��-�L �%Kp��^$�d���AX0;u����
�
��b��IE�"������� ͐ݽ]�S��3&;{|������]�y��N%T��T
h$G&'�L�J�J	�J�F�Nv\�W-�MIaB8P�Lf������9�k���C�ȇ,�%��]�Ԟǁ��NT�v��>V����`�7Y��z��3��ه]t�c�;�n]�	��˪�� �����-���)cZ먢���XU�(%kQ6'O:n�ڗ۞8� ��1FA$��)7'.����.?�%Ȕ�=�{�=Q�I�	1�K��6C(����ŭ�����7��7��1���ӣ����`�)Z���
����t�����u�|� ppp��k�о��r�!�ј���6�u�b6Gg�"��;�gw��Yܻ���(�+>:�s��ݵ�v��ԕ�����l�'�.K�}�sc����MRlH@?/뎫���/�eY~,��]VnY�V�.���w�^bDӠ�F��5��d@�2�����`?�1�����Y�is�H&�d³
5"�(,Z��=�b�=���qk�ZC�L����������ن�G�޲'��{�#±ZN�)��J&٘���E	�Ai�򎲶(Q0P���t��Zy���<{�G�;?y�����ǈ��/:�oU-��U���܀�+f�#�� �BD� n��,�MI�a�*,��*�d#��l*�
0BcИ�V+8*ϸs�.Y�QN ��s���}�޹�u E$3���[�wIV�%��.���k�R�&`P"�D�u�k��',�g)��=��2�C�6�(�H�R�,Ǟ{��(i��~l#G?��R��ہn��w�)]0��襱����w�)���|�� :�����]2�;�~��e�_ �n� :8q��&�gY"�њLD��VRZP�������~����O5��ڗʞ��T �S!2��ǰp]��9"@�D�Dۇl1S��6JK�.Q���j������*��_��W�
��3N����}����M�HZ��v��|�����Xmuõk�x���y�7�˓F��������c��%�n����#Ƥ��̍���_��Պ��������5�=�u]�컒rw�Qv<r�.d�>.��4��uY��(1���,�,��yX��e$��!��<Ϲ��Vg��9?Ƅ���1��Q�\;U[�shR���cd``!B�ȭ`��ߪT�Z��uR�h���!��A
��
-FC�IFÌ<�,����Yׁ:�[�����w-�sY?�ݧ�cAGr#�(�@+�tA)�'��I��̀I6b'+0Ab��AU	4o��!�E��C�%=7n� V�z��v�l�ݻ����v�"��[����/؝I� ��[[�����,D��� :3� ��(��ِ���ͦ�|!<�Gx��c+�O��g�����W_������������Z˝���|��I��u�ٽ��#�_A�֝�B�~���`$����2Fv&c|ԞԨ�<QD�V(�m�4!9��e��)v�'[��ܔw�������=w���q�6�J�-��u]?R����9u}E���("��>����Һ�r�J�bBD�1AX���ڷ~��|�G�	p��/|j_z�T��Jʳ��� �XDi�@o1(��l���2s1�25��o��h�n�pas��	�T�W�����~x��O��w��htH����]BsnJ��|�(��e�p�A��FG�"h�Ŝ�#j&X7��,����������c:9Z���j��ko�91X~�_���Q��|t��[�'�L�.{{���M>8�aS�L��`4(�Rt-k}�6_�R=z7���"��Is�����F��E�923    IDAT��a��}"S�3NΎp��DIUUH��T��\\t����b�ɠo��1k�f�b�YӬH)ט�>���]2� 	a�d�TPާ\����.;���+��L��>��3�R���f8,��&��K�JA-�2eHQ!U3 �į�d��k��פ.�4JR���Q��s��m���Q�^��Mb]pr�a�ƴ9c<�"c6?E��h4$<��8˚$#dMN&Z
��1��2)22�/���+��2�p���W��F��#��+��E݀@�0Z`�@���9�7w�B[�젅&�	�J�5-�Z"�Lu�~�Q�aA,-f�!W%�mL0����Ƃ*dM���iSsH����
�q���˺ϡ?�y��g������\Sw8�{��BF<BEv�y�+�\}v�`��w�l8b��ϲZrzr��{���w�ِ�%.�Zi�p�q���K��[����|t���������o~��vd�{��݆7n������Fh2�ϩ��9��x���P7'K��x������9 y�*L�b�W��jB�qYC�A,MI:qa���nQ��<UX|c�9�҄�D:�S��Aw�� X*��i!u]SU�:��֮��4Y!��1M�\hvی�D�w�k��U�v��#�������{}|_�XҳWkk-VX\+'���`�@{7'���$�r�L]=X�b0j��"E�Rx?�<��;����})�ɜ���2
DPA!�"&K
�պ��I,M� a�l�Ǘ��t~�B�X�ns������ZK�+T���d���]��%?��O0&��H�mp�rx��׾�7o^���!���|�������p��}����p�����l�6����stt�l�@J�.�Y���Ų�xmkC��z*�oG��Z��9���� �m�*�׻W�������E�:����-�~\y�m�AĔ5�ϧ����;>>��ÇX[���CYm03�g�����MfX�6��:|��V�*8B��hR��#ovM{��3'M�0���4y��ޟ��'L�Ӥmy� 	��᧿��B|�o-���1�=��2�����߈�����l;j#��<u��m�j���V�M��\[+�9E�>X琤�R�ܤ쉫+NOO�N���9�o�f>�o���,ţ|r_��`A& ����K���>���|�{�s��}��!U�� �@J����(P�	USR-�9;�����?��)�ߝn��ҟZW-rcȔ��Vܽ��Wy����وJ|��ort���`h��Z�)��1�N��he�-���˔�`������6ӿ[�- j�EB�J$JI�4D�xj���u��Z��mw㷿gte��-�\7�
�1$R��֦.�|���ϊ&�Ͷ3دh [N��t������0��	�bww�3V�eY󕯼��h,��yQ�Ri%�R���Nc=-���g�J�� Hݺ1����7��:�3�ݜ�v�g�  @)����i�dQ����Op��k�(<�/O��j�*�%�-�	$��>3��v��M�9�ވL 3� $쵀����i��������	����y?g-�p��#� M�`����F\I)���?�W�ݼ�c�蓎C����k+TU�{����ﰿ����s��9L}�� ����X�vv�������]�R�����C~��1<�X��˗Y]]mnސ�a�댛뺤(�MA����O.�>���	�/���S�p�9DS��pOR�}�c�puͤ��Z#��p���}PN/x��H����pt�ϣ��2���.����)i#�ik��*�ڢ�	B������nۻ�plx 
BZ�����5�W�:���h�r�lRQ��Cʲ����0����XWRW%Q��R�ѓ���<��K���O�8sp�ǃ���#u���6��IW�����Z]Bb]՝A������r���p#�p8D�U�4F��\< )Rx�18Sa���y��+�(�y���n�b>�#��T����.
?��צ��>d,Ǫm��£�D	��,���z������7^CĖ�9i�Y��*/*am�kCʣC޻�BL�B"�"J�$��V�ID?��#AY��{�%�b����q��W��M��O��n�٣�=J;"�P�#|P�.S�_��{���7��N4�*���I��c&�!*2�P��l-�鏮�]�+�څR�m�.|m���Сut���Ű�!�|A�9!�ɹӴ��/�n�Y�X,j[��ח���p���������`0�,k���)˒�����W�Z�����qB�}?��sc�'���O�������b�}9>����H�,f��%�ً�l����Xw[�H��^�BI8�� x��$	:ߐ	�#�5Rx����R�q���W^���+X[����-Y/�Ҷ<dooo׮��/�@��x��{{{L��N��-�89�t�C���5���Y���0n�m4�l�2���i��k'���,��l��$nM����i��^t�ߓ�	��{��ߦ�O9<�G)	ޒ�9�p̷~ɀ�!Hw���4�}C����Ǐ��ˊn�,�l<�p�5oj��`m�1%��Ԧ`:�������!��״���ԅk
��)�?a�M�ע}��������.yp����Ģ���7o������9���������
�Ǜ�� ,9:�FɈ^?�dIg��Dw�4��x��MP���Bx���.���oY]]����<xp?,^$S7�U���00�3¡U�	�]����h����Wōb�b|������|F9έd��t���s��w��}҉T1�%�T�\������B�����&/�>ZG��=�:bg�����l���y��"�s��%Dg�&>3�z�5�u5�G���Ѓ��Ak���ۚ<ː��L�@i��e{����Z'��_�)�_+<k�4M�� l�R!�h���0�
����d;cʲX\
-e����~Y��n��k����&�	���
����g�g��ё�L����F^:Q�z\:�+k�a�#�/�w���r�,�� ٠e���p�AVJ��ټ<e�Z��l4�[�;�B�׸z*�H�H��ш(�(˜$������������C66W���g���3�������e>�G�[��(��#����l�SI�0)k�t:�$�D�0[�Z[�ő\>:�ǡ��^J)ZT�S��|��Ok,�
=��]ݿ5B ![�k�̡4�������H�g�)2���Y_��=��pM"�r��^Gm�(B�A��£A�T�u֕8_amIY�p�0�g���P�9u-:�x��΢��8��찰[ �$/N�s�=<s5ݢ��t�Iӌ�h�$I������&:D#�GuH�1�4�H��a��h@��U[$Ƒj����>��t|�/���q�����	Y/���R�z)e�?��|�Z�
P1�&SY8��Ԥq��2�m�����X];ǅ�A���%���C2�IJ9?"�,YoH:ai�JŊ(�w�҂~��f�Dc*��7����(���7�@�����=��#���^��hfӊ�k{-�"���h%I҈HKr���(x�?	uW�H�k �"�_0l���4�n����Py!:ZBK%i3����5ݳc��l]Ҭ��)�<�\#fA�|l/�
���d7oE����@�mO2��������I�1�����a0��?�w���?�7�@J%�?U�����+�|GR�U�g�z�ϻ�����~r8焋��	�����^;V�=k�\�=����c1[.����v/�i�l
*�5����`D)f����cl�o��7��u�y�wl?z��!zK�0���!:R	���p|r�`�#Mz��c�8���Q�5EQ���z=&�IW��� Z�(Uw��{�@/�!�F<��(�$a}}���-z��P/�(._;�󷼂]F'Ϣ{�{�%;ۀ���t�a��q΄V��x	R;�ڰT�6+��O�kF�DhW.���]��7�� �X�\�?	�(_S�I<�U ��B8�j ʡ��69y1k��,���Y�5�O\��2H�(�)Yo�J"�bwߦv%��,�(jKE\�x�^x���M�$��
��ίG���H�\�t�˄βGH��)�����"��;��5E9eZ�C[Ζ� HQU�z>-B��#�'���k;6�'�
t�$��XW�d�d|�/~�S=�a��%ta�E�#._����\�r/"� �f��;h����R�,�x���'K&�}n�>J�X�or���Aµ�����(&������dDD$:
h��p���\Acp��eLxk�!�z��by��z�E�vQ�=+�m�s���R\�����ͭ�W�u�֓$a���Ÿ)�H�p��.z��M{��\ӑpg�ݟ�tY�sJ);���xZ)�9:<A*����ß�ٿ���&k�k8�y����|�����y.�2�x\���NƫZ��*��y/�/�{<�cC�$�H�{�Cs������ܾw�\�]}T;����27�)���KE����4���b��d��T3F�>[�׈#���ڵ+�e���;�*��K�$I@h��G'Gd��,���$I�|̙#�t�܎%��
MܗpMK���-��$���b�z=��{KQ��,�����E���#}X[���^z��Wd�\5��%΅8*c�MF����~��qO/<��+A����f�ǟ�N!��E�bm��AZ����Y%]�^`�����Bx��g,x���Z���эi�j�oQ!@i�w5:��y>�xC��A`a<�~�˗�r��u��~��*��)��y��:!�����9�PQD�#Ԓ�H)�ܕM��7|)C0��iLU��"CHRTd��ȃMt�/,Z��s��N����炝H/I�.��zNGr��o�����h��G�$��`��/��*?����À&'}t���T�Li��V�R�,���S	�e6�p��ۤ����&�%��fl��1�%L��G������;4�}S<c �|>�4��`d�MXT�3���`��8��>��ܙ4����	�'�
��3�罳�-����P����8f���M]��g���B�ݽp:�m�����p����$�e����U�慗^������޿����E����l����'T�%k�ON���f�p��o���ّ���������8�� ���|B|\����y��&�m��l�p
-�
0��:�o':J��)5ei��=�ш^���ã=�6���~HQ�Y]q|b�N�E�x|�(.�
{>�vm���SJ��=��RW�i1ĝ�_�<�b1�ڬ-�<�ǎA�HR,��Hwj�e��PB�z^���/�����f���l�c���
(h�w�E��ؐ�!�,P+�v#�@���x� �g�>�pq�R�A�~4�_���_��x����	��U���(=B��Ƙ
c+�(%I�"�����-U��-G�$�X<��^�|6�Z�"M��DQ��|�#U�4MYYY�r�[^T���yM��*�D��'ME	TEG�B@)��u�#��7� )ΦAJ�Ғ���Ee1u]1�N��dYFU5|�S��pm�?�L��o�z�	��H�{=I#tB:��b�!N��g)�����c�jfv(���o�k��X[���
��#Bb�R�q!=RA�UH7�X�� ),G����M�^����*����Wz��x�T�y�uQhѱ<ϙN��u�Vqb�Ž�H��w���{\�pCגn��)��Ej
��s�2��}m0X�\b�����9��.E�U�.[��������i��M�|ip�m�T�<���SǱJ��������o��K/����XҊ���ƍ�z=����r�
����]�u]+))CI���[�[o��%��/d<W�W�W"�8a�qRD�*�,�cP���^�����G�u]s��e��~C`?�����4M?���J��O���2qj=#QAҴ�wtF
�����]h��Q�h4"N4U9�~�cv�k�����~IQ�qƲ��M�Fx'������3��9���\<�۷owh��񄕕������_kݥ3�E_Pg��7��9ٴ��ޓei�bmN�)t-;��0!'���!�x����*&�6���>��g.�s�>lϣo#�AW�5)*єEN&EG�|��V��!��w U��-�=���H���a4�ĺ�JP�K����>\���eN�X[gZ�@QU5UU�kT,�O�j���>�R�����.r"E����Ue���e�
��������}�����+_y9�9ͥ����
��/��n�]��BX`���c��L���2����3T��~kmC���������X�<���a�W�K�ʃWbʺ�zE������c�X��:!JRfSà��&�	i��%	��q8�^�kV��^3�`��]+e���eN:L��qrN/Yc��}���?!����_�7ڢ�'�B1�b��.8hqc
�kx�H9VVW�(�g�4^�?R�4ee�����:�'3��)�+����g�Bт�!�[�����,K⸇֊�*O)w�E�֚���Ά(̹a^L���ڊ%���`0 `41��-W��W�!�i0���NY���c�$ass�[�lnn�2ڠ,K�޽K�$lmm���#��9�� �����ϟ���<�y����w����Ue:�<����>��6�����R3��.���(k!���j\��[o�u�c�_�/��x1l��.rRJ��!��{!�Ctj�g=����p���*eYvR�4�U��SѐjC=�lo��@D][��7d}}��QG���G��,u]��:
�#��xb��H�&��7����t��YAQZ���7���[ᵫ̎ /%R��Izy���B���e�}k�ܒ����/�h;v�N�[~�?No'�4MI���F9�������v�פ���@h�FQ�Pck�
��BL)�����q���C���gg��'���/֗9o��k�����V.��p|<���)%�Y�|>'�Ť:�,g�\�φ�c��*7�%*��%���.�э��sM1�	|�Ó�o��,��g8Ҵ�Z�"beu��h��|ʠ��7G���(퉵���3�X����h-�g'���?��0�!R��Sa=�C$<�/r��98xȍ7�<_ya�A�`�D��Q��	��#/
��#/B������67���!/K�
��F*�$UQT��{�a4X�_��&�^�m���t����;�YƬ�hP��e��cNM+��L����;w�<\����j�vk���v�P*�R������0Y���z�M��������
��x̵k�XYY����{��Q_�����׿NY�ܽ�����,���{ܾ}��lֵ��c�w�9��\8�R�ⱃ���g=>��#����(�9'�t���>�Z�\~��ڶ��<���ڂ�I\��c�p=��cyH/�v`}/jՎ�l�����q��9VW *lUr��<�WPy@��-�4%�"VWG� s6�6��v����z����!�������X�"��-a�Cv\k	�ϬtR*�q��vZ�;��v��E���,ӳZ��X����+�jS+I�$D͝`�A���l��V�'��h�Pm��2V�p�!N���uЃ7�0��]-#�tqv>��}�t�d�?��%%��-m��f���6�Xou��s@���&��3��L��j�v�U��B(�X��u
![���"�T��M|��Zy�%���p&��,�B�H�n#�~�CE�աɋ�8θp�*k�[���*
����
c
L='�)�������_{�e���]��<P�Q@[#�p8R*��J�DxI"�ق�b�g>+y����%��ӿ~!�H��TL*��(ͨJͬ�QQD�E(o�r�:_{�޽q���Cjc���'%�� qD����~�+|���y��5����c�ݽ�/�s�ܹ��GO?�˭�v�߷T��(�⮋����K�\өq�u}rr�xr@�e"�)q�q��Z�|>i�C�1��x���Q������p���z�%;��Zs��9��kkkݜ����ŋy�׸t���ܥ�-k̋P�~��_%���w�yYS[h+:�Ҍ��Ka��3!�!����e������+��@��{JJ�Fz�!�    IDAT�{�kZh�����c��<�>eY�]��J�i� ���>
^bNڮ���dx#�d逵�67G�R��!�uf2p����F��3�i����e}�!i�����pttDY�$IF�$Ե�"�Zr��-Ue����C��Xۺ;�SEA�&��hbA\>Mv���RH6"�� g�zZ�x��
=����E9 �M)�w�)�C[�k�@�7ކ�)��)���v��E�v��:�v��`Q�dԠ{B@��=X���<u(���R���EԡގP.�S3 䂪�Y_�`}e��ׯ�#RM��!�7{ё�E���+�ٴ�'d(R�u�s`}�ݮ��6"�.�~���"k+*Sb�'�R�b���׿�������g�lz�|>�N�x�E���	�ϭ��g|�O@I&������ܹs'x�	���x�w
SC�N*� c+�g�d�`�;�X6��Ylr~m�ee�ޅ�T��NҌ�L�����4����.���}����<z�<�69��A���k���:���&�뛬�mP�5E1gw������?�1�*B������D��A5)0����ϝ�E�ϟ�d�t:%�SVWW��stt�TS;t$I�^��
 ��1�O(�^�h�JU$qF�FL'��N����s��9^x�&�	{{{L�S�1dY��/��w���R����|pg��/�e�yAkVVV��w�y��n9�a��B΄RR���������������/d<�zw�Z���.Fh'b�E)^
�&����1g�7�2����jUP�;���YV�N����>���.L���*[[�����)�6�p�2�M����	�X�,�ܔ
7[QT�e��G���<x��������'�s�$aee)%��PH���[�!���W�D����}ʘ:���E\���!t��8�����X�7y���BȝQ�6�^�cl~_iI�e�#}(V��(a2�
'�Kdѫ`� !��#}c�,�`�9����ؠ�E"t��-Ri��o��A�#E���g�������O<�X6ŞpOR���"HVV���7�䅫W��S�,[��pO�:�d�T����ĲD��
)u���'�"�~�l��l8�A�{����F�1��i6o���ˊ�����]�_;��)��/w���<|p����S��#��6YY���7�/}�Ud/a:=$M��}�������Q�BH��Y0zd��R�%��	�	�h����1DB�瞻w-�l�Qo����YJiJF�b��T���jDl1N�Im=�2�G+���-._�y�c�y>&���qJ6�&}��h���j
��>�����׼��;��:j���S5��Bt
�6�m���pQ��-�~���z!TJS��$I1��(Jf�)�露���{TU�����\c�CɈ��sD��L�ۖ|��Qy�wԓ6`8���	��.{��
R�e��W(���7o��H���q��^�=
!��H%Ơ��
����2���k���DJh�X0�}��]��=�}�����$鐦��i��5>i{7�nИw����H��b��367.p��UVeuL]嬯�S����f�&����Ƶ=�1��U�(q3�����`g��,���*���7��q�"[v�7�4��c�E����/��j�Ek��i(w�vN>��h��U6��SzM�P.dAl!���@��+�� �B����}ֻ��N_*B[�
"I,.\���9�R!�-w%q"�����k}#
���e��G�!�
���]?�}�g7�yE����˺�Ը\2��ڵk|�+�p��y�j�mK8��L��k�m��k��N�nz���m��YxHʈU�E�DIL�H�>�����E�aHe9�������W.l���`�5׮_a2�g:>�*J��D:c�_ޡ�����X�(�G���������h)0U��B��t:�,k�h~�d<g���$JgX#��!��~�w��Z��n�z���&�����u�ԜL��Uh#��"d
u����c�pD:ec}�nUR�S0A|��2��r2�b�GE1eY����O~�c~���SU����i��\���e��5a.˒�|��w��҂{mm�_|��xʝ;w ������A�M��$I�1O��ʾ(J�
?��666�R0��h��x����8fss�8�I8��=���tH�ݻG�\�~�<��ƍܸq��vm�]���1���766��o��eǿ��\E_m���v�:@�@�RI�r"���=�[H����8[�곎���}��]�:�eMU��<��y��@r|R3��p�,;�����\�r���5��)���[��r�w��9���ܽ����}N��R��X]]Ek���.'''$I�e����J4����*���->����=^���O>���w�����+�˿п����Z�F:�
�X(�������</B�֫���@4�7G@��V�L��;�s{f�p�$����*��ƣ�`�ӝ�%.��is�������Q# ��g48T����
_׃��3�c{{�|:Ai�|�\W�i)�.X	}�l���i�K�M^P�j!���DЅ'1^���ț�v��SCu�g���w皮m�O]��p�&/����?o�ƛ�s���m���>���Ջ\ؼB��ump6(r��)�uă!��~����o�����G��\;�xf�`:�3�嘍!�d{g��}��T��e���H��*���)^&��7޻��`�H������?���gQ�B+*�8>s��
Q�����xj�+�tD�`�lBR;�`o�����;��m���YY��e�uIU���no��`��v�B78O���H��TY�M'�/��� �K���8Nq�5�^AQ,l��:�&M-i1:+�V���y�3l�ᬵ$I�����C��@����=N�˂��u�(���9�Yjk�D�&;�3k;E��я���S�������H�sBi/�PBJi�.<8E�mbiE���K)�!b��z�4-s,�g<O{7��<�D���;�,KI{0��u�����F}�^�ʵ�3�N�˒���]8O������׿�-{G�$�ek뛬��1��893�Y[�h���[�Y���K�e�/�B[�"2/P�Ӧ��b!��=�����}�Gl=�
��m�h��"؄���{iz�$�eKhLӚ�h�q(!2�x�bmMU�H)�W��s�7�7m��\�E݈�G�%�?�aX�-��|Z���'��%tԇeN���oݺ���#�8��s��Y�^T�Y�	�7�\
%�:>p`A
�p ��&Dg)�2'�ׇ֤i�S�e�d2�,�ywjۄ�r��4�-P"�ރ�TE����M���6FԦ+��xop�RW)��u�DhE]��������.����gS�xE�:ؓEX8V���CƓ�y�P8g"�������W��[>�����VV�ܾͭ[��̦H����3�Lx�h�������T6�c#"G��CV��,��	4��䓒[�n������?�Z���j�zm�"$������{�庵ܷ�a�h��s�$a6����o�����$	�����j���eMk��q�z�eeYrtt�|>��_�Z�I�0:�s2�t����ۦ�lmmq2S�y�w:88`ww�?��?������g?����.���B:�]�p+�l��/�?���E_m�L����9Q�8V�>ʍ���F��DG�<�i�cpQ�	��e����`�P���sDh�Z'I�U���N#�	 Q*A�cBJ���j����Rtxd8�_^�M��y�wv�ȁ���d����ܻY��"�J�[�_cw�psJ��q�ҋ\�t�G0�?�dg����M67C+���ܻw#������k��1�s|r���Z��"�S�ӥ��S��Y�m�kreCFr�1P�_���&Uh[C�C��d�MVd��|H}BӋe��Z1O+��OA� C&��|�><yq��ƺ���I< R�T�GD�,`j��b�^�#6�]ccm�)��cU��4R%���c�$l�X!B¡���%�[ba�eN9�G�>��H�^<'�%B���S(J!�¢�EKA�<G'cD�%C&�l0D�����-�Z��Y�׶ЯT�����H�P��v�pB`e�P���H!Hc�)r�|LgX;d|,�	����9��l���A����`��B� pr"B�^���+����r�zN;FIƴ8��H�r�2#B \N,���)uY���^�э�Z���M��'�~�uQz���s�QMP�` $��}~��cNv��Ͼ�o~����$!���%Η8�k�7�y������_���Q��}�V�z�kN�czf��dʃ_�7���g?��ܕ�B��З�K�Jcs�4�H� I2�x�w���=���>'''�'B@�G_D������� �qK7�AtH���:�^Hp1r�����#}�-��`��&ZW7�8,��eG�,I�P� ���ׂ���4�ac�!<��
Q�'Ix%��$�Mf�	u=��_AG�a6-H� ��)�+�p
8B��`�'�F+8�u����35�Tp�Σ�$f6�09�Q"���P�N&��"�bp���\8w��sx`0u J��yI�qIQ3!R#�Y�)2� E��;?N�'�5����_���я~�I�޿_���E_��;m�y!�x�W�[��y��Y��
�۟����a}-��JRX�����w��������"J��C�:��k�X0�������Ehlmm�ꫯrt����i�t:����loo3���hD�$lll0��L&݃��W��z���e,�-O0�?�W��/H{����AkL0�n=c���X��$���U.]�ĵ+�Q*ؑ@���������{�j⤼k�=��FKh�0u@�A%8')�c<eY!�"K��C����A7f-�8d��U�)���p��s�a��G�P ��� u
T"I����Hc� �h�k(~]��@zZO@���X,"�'�8L���ru�{�N��ZŌ�#և#�sN�w(�YE�k󳞌�2�rHx�Rz�j��;7����o8�"Q�%���5Ζ�C*�������������%����Uf�O��O�͛�(����n_�����K�c�R�RAY8�u�S圌UY�_��� ?���
\�5v�D�T�M��+���Ռ�*��>)^��-Fh�6�[�:�D* �
�-��V�I�`�
g�BL�1E9�*U]�l�=)4Λ`g�O;�V��F���c�ܹ�p8ll^���
NNN8::��իH	q��c�ֲ�xo�L���P�U������Z�S����0���oZ�WF�QE�M��':�_�/�x��#��JL�ｗކ�+*��v�mզOg�C�k�i]z�rw�Σ�Y*�"�x|���3���ˬ��o\��>��`u��x��ct�cw����;��Q�
V���[k+\�|���-�s������n��޶��� ��a5ݴ!����=�W�l�v�ǭU���j	���������b#L�j����A4-��[H8O��|d����ۺ���E9���T�	�m�k
i��Y[nՋ�M��R�(�J!��?0���d���>��P�B���I��R�$��X�	�����I�/]��ڧ޼gc�����6�]�h���A4���*1¢��a�����@^�������2�8��
��"��rw�*X4"��� \�
!BKLـ�{B��V!��Mr����{���/��M�^��)����ȝ�ߡ͚������O�̇+��"dDGo���|p��7�)BJ�g���]���������h�XOY�sgkL-�#�3��wnq�w�Z�e}�S���J$D�	�����{�K�8�RD*9��Ԧ��΃@u����A�-=�m�89��!�2�V��'�^�w��8��K��ҋ(5U�1�ƒ	kPJ൦��࣮J�8B)��hN][��5��'��TU�3��P��JE�klm�u�q5���AG�Z��f2ws����$x���EenQ2�ʕ+!�c���l�e��r>X"9�!�C)���D����U�EZ{]
YW��*�s���e�VE���3��\��{v���HN�"M���������o8?�����V�׸�R
Q�������.��qtt�W(-��bv�<���f3����`����k�G�8�"��޽��Qh�dY����Y�[O"з����;����4?��?a�Ҏ�3RH)�|������;���>B�< �q�R�5'�)�*q�P�-n�D	2��Ea��z��������=�$j+�k�����}*k�+�s0诒d}��*np��j7$SHLT�E�fߟr���=,l~�X2�>���$�)�Z���DR!��U5UQa�G�4��p��iS�36l�w8b�p�" *a��8A"p$�uH,J���օbNhjkR��y�7���]���g�c��e:>��WDk��Z�|N�,C�Z�6�u�,�����!&��:��U𜌢Z�]�0t�`"��KZ�4E�R��Q�,�b�>j��Z��mv���Jΰ��ƹ(�J)��!�E��`	~�����2�rh���P�8��0��\й,<�8�i�"�u��WW��RjSrr�d@7��$�J"EP𛺤ȃ�6�����c����4~�g=:RX[c]��H5�3�XF8�I�OӔ��5z���T���u�]�v�S��(�Nk�ׯ_g8\��������ˠ_�sNHD^?r�?���s��]�_�/��X1lxo����ށw8����[ŧ���0�^����mW�4��n����$Iё�*s�}��e��䐣������>�"1V����!��`����d�ݻ����X���#N���'�F�΋��r�����{97��� �g�E���S/4K�x�����޷��l|��llm���m6�%�f��W�d2~�Vo]�����1��cY�eY6�����lk�[/qޅD����N�m^�0�����9�{�N(+H��N1UAU���\Y?���*[�xW1�3�}�No,^�<�gi�x����Q9��:���$�ܮ]�ֹu^z�%F�!�*�{���7?@��Jǚ4ӤYL�hL�֠T[ny�M�ƅ��&� pE��;�u��!����|�B�Ƃ�2���X#�2���Ο?O����p�i�R=��S���G�C[�Ra���!�$R1+�Оs�x���\ݕ���uU��yn�nh���K���y������siKyP�1�k$�������Q,��L`G�"�r�k?$�!d#l*�X��R;��}�rY`���8g�Lf8<Q��T���4�#޷Tp�P�s�*u�J~��!�Bk�X1�0Gp��a��$q���.%G���tʅ�h�%�akѴ�ei���̦ަln��_&�2���!�E/�{����[�ȸ:��ϻZ���i��U�E�H�z|����g5�nˈXˇ;��O�֗T�H��)�Ȉ(N0u��7GQNy��>��y�/����pm���&��)����bw�$�$qȷ}�hֲ�x��js�����c�ݻ���4Mê�1m�ܜsO}�/?��|Z�H_;�{��EkW�9����u6ϥ>dg�7n|Н�`$l���T��1e���æ�rݤi��p��o4^�vUz�ex��B{L%D� �$q�f��H1B
� "�z��mq��6�G�ń��-D���AC�5*8k��c���<]|�����PT�._y���/����&��	o���<|EN]�И����*��d$֡ �B�����(��Ix0��z���Fk����2��`�(����VV�HӬSOJ�9],|�����є�ߴd֖�F0�.����f�u�>ȶI�-EE�s���R���˧�r=��tu���,��B��s8�R^��HJ���=PJSzYڨ���D�t$��l�1�,]�U�aU��Z�bzα<��=,
��p�J���$�2�@�8jP��؎"��I�9�Y&��2���P�7]&Ѫ���P���2M�\eQ���O�����    IDAT���Ԇ�BE�^�Q[��d�ݣ�h���!�-�s�����k���sOe�ɋ���Do>�˷�*y�u�����������]�IQ����E-�wz7�`]&�����~]V.�����KHIk8�M)!����	�]o=BJ��y���7���ܿ��/_�W^�ҕk�C�
�#�*��!!�Uak��d��考�Cd�:i=[ې�����8>>fuu��ܵ(�2b����Z����(X��I�0���9�Ej���H����[��j泄,��d_ꪤ2QST+�dY��/6~��T�Y��l<�hb�N�f�=�I����� �Y�G�*�:�?����tF�KA:<c����8PY��4Ր̽���3�_�-{�M��i�D�pT��NJk��u.\�ʅ�5�Iƃ�:�����fK�$Ǚ�f��g�%#"�2kA
A�
��閙���6#-���as(�&� X���K�q_�L��������\�P�����Wsw35�_��T�zEJ�k���8=;f<��i	;��%�=$&��F�L!���Llq�������e8��*\�K�
��z��(�uU�F�����Fߎh_��!MB3g��"c�R�&��_��s�h��$�H��_Wh��z9�i%ƾ� ��s�#��T��wl�*Ꝺ6�i|`��o8}���"6-o�M�GB�zs����(W�}���ZKD8x�o��ggԭ�e%#14Ik7J[����A����F4��$;^�������%��7�&R/J�+�TiL��{�0�r�F�F�	�˪�����j8xu����'��ƛ��h}��MRoÙ���b58������E��_����gj�k���sE���q�j��TDt8��CY�޽�_�1I�(�0 ��]���Ʉ"MS�J��Ņ�('g�{p�������aww��tJhjvv��7Xq�JY��'�X��O��h8::�6nݺ�b����:mF����6F��1}���Ί��<}�^��8ŤX��R���p���,+R�C]z�y���6k�5,b��?ˌMчˑR1���0����!�u]����x�99=b�\�\�h���^)kOU���h4aR�t�4��Q�'��WH�iGμ��6J\>Ƹ���>��Yk�rK�;��cLPW�D/��5!:GU��Fr���O�0*uS��y�&���ɹ���Ȓ²�9==��|I�-(AK�۩"dYF�4����K�}{�y6Zs���3X�D^"aP�Fw[qb#�"�C$��/�����|>���ʑ�%������R��鴏���$����1�k�HB���Ɛ���7�xc��Iz�I*� �@Q��k]�Ջ�U��a1G1��������O[����.i�����3�l�b��Nz�Q+����ELr�TB��E��X�{^�=�T�D�\�9˻�ڐ8B��>��!G�f +�x��o��?����ۿ�?���NE6u ���0���$����A�AU��9�I<��ݻ߾P��}-�LN��i�&�� 0b��(���0�M� mp�O�1��*:C����buI�n̼��X�sB�r)�wi0%�UD��-�FŚX.�X�	wr>������L&�f3��������H�h�4�r1g�8g�� ��Î�S���y�Z=ٻ�`�&��S���v1����]���C�`�4��q��}����/_����p��o��S�l������*�������w��DQ�u:�&b�a{{���{���?����px�"˱VX�k�Rb`�Z��Y�	��-f)u��Q�Ν�����VG�"�G5R�%*�&6�U�x:��+><���o0��&����������K��xL�˧}���N"��I�[5/�u�|4�mEȲ�,P9�3n��g~�Bb�Ν�L�...cs��f�Z`D��g���E���)�#vw����,��`�Y�
����`�� ks�/P��1_&�k-����] &�IOXH��*��ϵ�0s�>�<�=�z����8��2x!� ����E&[�lmj����`u���צ������z�]thX�}'ǚ���.=�>$bmR��\F/��ϡS万`��@�o"�vi��:��E3���];_v⾲y��V7u�s4u�K���S�����O�ۿɽ{��w�GY,E���9e]��#�|����;;ЄN^-I�9�R� e���pĨm�Vڬ�e���ֶ���_ݥ��I~j{�K�mmm1�88�K��0�Z-�:�A��՝|�Q�8�IفT�8	�ߔ��������m�?\��bϞ�5Fc��IPE��FU�����d}q��i��j��{?,T��cJO �����b�����|b�O��\-�,P]2���h\���2�,'�i�1�TAhj|]��e"X�����^F!E�5k��!fo���9��2�1|ݘ���y��H��6�(��qy��M�����> y��U���S>��C�5�Q�%��Q戡�)rG�Y|������c3�s9M8??������Z椴Ѡ--I�T'�:u�J�g	[�����1�0�&�'pn\akmH�s��6��1���S��Ӫi����݄�\�-�g��}dk���[��1r���w?z�Ç��u���� ��˳�^�&'��� ���򐲊�z�~rNc�����*ߪ��~�"��h����E���37�T=����>'��~��V����Sr�t�o3z9Z�QP]a�z���?���7�q�Ǿ����Z��^u�_�UU��kqy�G��>�{�d#v�n2۾�[o�`]��~��_qrz�[o����{+�R��I���J}�&����4Ep���R��)�g-�ṷ���2��s�dY����܄
�2�)�O���d��D6���,��C��*D�چ?�{��o_}�����}��Y��Aϐ���i"Ĩ���vn��:���U��u8�LY�E�J�YBS��K5m�.����^�ΰۊ5��MZ�t+-'�q�Ybh�c:�my�4z,I��� U"�敽�#��(�X!AlZ�s��鰜���fD�e�����ڶa3�U�b��5'ƥjHqX��E0Zy\"��N!rz��s���ɸH��1�!�����Ua<����$��hR��������YT�Ծ�	5j�@����l�ɇ�)�kmJ���{@c-�Cr؞ކ�޿���m�5���|�bQc�8�������F
5�"�$��S��)'G'���;����T�yn������	���&�-b��V+Bp6�(�LFc\fPm���Ū�,kn��:ǯ�����T8m�g�=JQ�֑e0�ʠ�;�*�r=m�^���������Ē��6�k���y�?�%�9���_e��ĸv´K�>����f��G�߯/-���I�Ŏ*�Q{1�/�s.�	-ԧ���tZP;y�""qMk4�VLg����������&U+��	�4MCY�}֤s�D��h�!/:�t�eh�����,F,��͕�o��:�ҝ��c�*���g-�Q��朝�%�WǛ�T�*A|1��h�yc�v9���GGx��}#�\�>1�bLH��h�4���u������������t��~�����j��N����z �1��)�D?�^h�bM��9�X��7�/���:�V�t�&�ۑ@;�в��g|F��q��k��"��k,�,�9����(OSG���]�G�<��6Q7t���Ʉ��m��xRP. ʍ�=�g��i|�3��nN��'�
ʺ��!�Fd�4�ȊU����prVS5���і3�f�,s��`]�E%�{n��i��^��N���t�~
-���g��^�|�^�=E�k�8g:�2�LZ'�����rNӔT�_'���l���=f�m���lIU՜��pq���R���D�!��4�r�����������X��Y�-��ç>z��iˡC��1v�i���4���9|O�0�����A�n�fi�2�}������`K�Mj������u��f�����Nx�i����K�/fݤ�j1�ĸ�uϲ�Xe�8$��$Bu����+.3�
��F�]�nȍ0�nq�`��I)z��ɰ�`�����6��7i;��Ј0�'};w�u�	x��|_�d	���9182;�����������{rxx���uT��i�U��\��D�ЪV�������1a_�wƞ��+K(\��[pѪS�(�����M���a<O��*:|"����%�*Gz��cl�N�`p�]H�U��~9�`�z]UM4�1U;~@Y�pN/��_�:g�q���'���w>��F��j@H���
�s�b��T>2��:�@Gm�e��J*.���`gk�ӣcV��q��֘���"����HSVI�c�3*�c�mHU��boo��(�ǣ��D9:>��	H����s����F�[�Qf[�:���u���dY{�����(�:�W���6a`��1W��l|�*���o���os��>��}��Pΰ�����;�ܿI����9��X��Y.眜�2�� ��l<b2as����a1_�������8:>e4�0�n���o�Z��֭���)׍��#�tU�=M�^��I�E�L���c#��'miQX/�X����:F��=à]_��+W�b6+�t��^/���c����\2B i|���`����j����A�n�~�����9��sv����C��n���K���9;;�В�'j�%�D���y��S���o3AI���x�����4M_`ש/ucbwm��L�˅�.���S���|ʃ���J�7����W�"j����y��7�J����1}"��N_�@�c�&��VET:2��e�(��һ�s��%�rլ�{��,6�;�iYόe8��n�?��4mg�!jr��t�i�:�����d��aV���_Ԇ�Ʈ��v�P.��e��y�q��E�����m+}2$"!�7��y�=�2�7�N4���<��s^y啄��}�|�5����8?9�p�î�|<��<�f�&����ck�1*�����4JR���l�b^��H&�c����2�Hd�loo3���&T�S̏s�z\g10m;��t?k�d� &�����c"pzzʧ�~ʍ�XqL�[��H��튐�U��PWy>�(<���V�"�!2�looc2a�UY�������>����nJ��bLh��q�i�ez#M�m3T,b��ω����˟�*R�FV�z��KP7h7һO�Fq��W����ٝWM�0x��� �@@/E��	������7M�#p��=�������������G4��r�r��^���s�>���N�_������HQ��������`B�������h����C��`��Y��������u����KwOuϠ�TU�0��+�DL�2޻q���%�M$��Tc�Ce$~*�֫�m_T�Jl*�,N_zG �[�jT-TԈؐ�k'�_�+һ_��=�#g"������Lb���iA������1��i���V�4����`Z�!��EZ�-�i$l+<����Cl;��s�i<�����0�ڞ�:Ƙc_Rvx]_�6a�ԆЦA5�DIn������GTָ�>�m�:ӟ�l6��A?�����W8#_R��0Z㌧Y�m����R�:��l�+�^��믃��?���^P�D�z|r�r���"��S�RMkgyb��s�a�x;��)n��9~�hf��ެ�E�,IJ'�iSD��'Y�UUE��d�`>_��_��������wf4��������8�Q�5�ɹ�w�����IJu`~v���G�D��Ŋ���G4��9��>�7�S:,T�Oc\b;��m`�b��^�]֞'�M��TXs�B?�4�}`�Tn�E����v�-o��"�_y�p��uI#>B�4�����e��@ދ�]�c�i����c.V+2W���~�F-gN�4�[5%#�|4�����ƍ�N[g�:N&#)-��#������>h"�6.��Y��ݏè�p��uR��Q��k){Ʋi��9F���};�Y�*ĸ2bVx]a`|�c
.^����;c�髍ё�ob�@FD4���}O���������s�����e[�aL�'��֮HumD�����������P�
=ۼD�>�m�vm��k��6gb/���0�������P�4���q�����4D|c͢�^�$ ��x��J&����{<M�e����9�W?�Ï>����������-vvvx���.W������!���Lfۨ"�\�|������Sמ��)}�^��1;�3�����6\RGY.�V���b���?�=.�$�!���u�,��t���	=�1����jU�8��jŗw��T%��2��5��[os���+|��(V�U?�؞mQd#&ň��4e���!�G'����Z��1�ęƦ�����W������v����Y�y�a���!�}��9{�J'":`���G5tYߒn��#�L�١|d�+�y�o�X�c>��'�(���N��F\{���ØV�CM��� &K�٘�2�/�X!�`4�����KCţ˰c>���.Ҽ.�3���1}�҆�	�����᲌�Y�Tvs����JU��>��\.�hGp�����39}۾�y�b�oauo��is��MY1N3�^�G2I��I�H�>���(O��^N�_��i�Ä́(�j��s@]=���YF>m��2�3���A�e��TU�)��G�Sƹ��(�\O�k"RU����]w�Wo�}��0v��h�����Rc���]�mM�*�q�MlFn�(7h\����qt�«#�r|P�
�qN�8����Ҁb��U���~�����U����|A�q�:6�9yh�����{_B11Gp�Lw���8qT͈�S��E�qc���?d<��ζ�|�޻���T��?���l���>O�ٚ�(k����(˒y]�}s�7f7���+|���|��g���<�����u������P�S�m�'_��ݏ���)u��{�����l�'���Ԉ����`" S�QĸD�'%�ɩM���9���޾�b^bl����P����)�{�67��g���/������?��r����9���|��f�n�����C&���~��� 	�b���Bye�&Lw0�Ġ��^��j�B�*�Dm5E�::������r{=-��I����Ϛ�j����^���a�4��t�|�
�[�/ɰhm��z����N� ������e7�=1�Ք8M�\r�6�Ԛ.sqUA1Q圭��O��l�E�N!\{���؀����Q��^i��
W�+B�&5��(+��?<Y�c���5�pb�pNaGԥ�.V�Te�J�d�f�pqv�a;֋Cʪ5�D�����m9�wo��G��[i���5�^����0�Ƭb�=Lt"��J`�R:�k8r �MD�W�� &�J'������*��)�#9E��m8| (HletB�rhq��I��E |�  ��vM8A��)nI�Gy֓z&,b@0D ��(1᪌ &i������t�0*����JN�>�ͷ朊}��w͆�䄏[߇]Z$qߥAŵ*[[[�����l6��4�����bӓ$�q��9�����e@r���{�������^����o����O(lRI0��j����N���M���/�h�hS|3��}?�N���_������6�޾�̓vv��~倽�'''|�ŗ	�8��n���::�)�^�L�4�#��B�A�}*ˈ`�
�v�=�ھ~�\�z9��}?|���~/;+�����q��5|i����-��>F%S�L�#b�)3�\,��ݴg'g�&�Q�h8#���D����3�` I��|҃+(H���Hh�Xc��Φ�G���9�˨����YKh&Wo�}v̀k�c�f��+�0��.5\.�]
$E�������FWfɚT�P�+�8�ڀq	�d�������,P��'N��4Q�t��N�a��x�R��� �Ι��ޣ��d�P�ȇ�����{�p��~+]癴�xu�`2\6�co͸u�^y�������{�����!�}�E��N
��d&�t��A�d�_�>:,n�/��۫R�y��4�b����=��o���%�A�    IDAT�G���p_WM>��3���|�rV�
I�Ay�X��Y҇c,J��'z��
^\��4MC�U����5a�|�_5x���=jCR���>+uyu����w�L������=iR2<����{�o�IOAT�(�QSˊ�k8�k�6�3;}���L'"���1���RŘˎP7x<�����FD#N��ƚ�K$4X�����W5�b���V5h��J���	K2_��^��^ds�VZ|��B�k��+�S�;B�QR䍎�?����l�����Z���@�^��f��"3�Pb�a�[vg�>��9��S�~�Ï_!�s'�A���I���X��>˲��t�R���;��w~����6�u�i�b�[Lc�m��@S�d�e������������*�5Tu�u��M��0}�M8�C�[z?�DIҜ�>6k-2��8�kO]�,�Kʲd:M����ϗw?㓏���Ç�:`M�1	C:_.����h4��H��D1��SʦS'H�^>j�V}t�9m��c�������t�ۢH��j�(��0E����U��{��l�yl����R�o8��!h1�%� ��K��|L���]�g����hM.Q� b�1�1��nVI¦ӇHO.��fEQ"F����$j�5cHd�⒟��ӈ�R���*�}�>� ݂t7_��&>f��!JΡ F����I_,�JJ��$�ISVT���D7@��`���|JrGѐecn����ɛo�f6��fNS��f�Gºk��~7��4�fg�~���rJ�k�,�h|�Ӕι6�k������.��$1��NP]y@�l����F#[d�A ��
[����N'hU�%�O�'F�?'���o��c$�L�d��9*�pZ$U�Z���>������!��Ox���s��O����9>�G�elMv��a$'�G,V�t����,<h��BL�Fg����X0$^�.�����3d��{�����[�Ӕ]�y��e{������w�.ߟ:p���w��o���Qc���(��]۟�=���C'Nѐa�c��D�-��qc�ߤ"O�{rz��qs�i��C�$��a4���
���k�T$K`n�o`�.W j���ҿ�H_��cΣ��7!`���S1��	m�"�fkUi��#bɊ��h��%,"4gyR/(Ya0�`3G�a���o��7�џ��;��Qk
g�)���y��6�B�v��"��6#˛i��:w���܍I������Z��f��k�1�N�Ӕ5>(��+O��XuT���sm1����6������՜�B�S�f������d�5��R��H�_�e����$|��]V����|���x��Œ�������������x�>xL���Y1����y���̗+���4��ڂ0�ku3�Dvxͧi�+qQ��k���cCxA��x�^^���Q���?��5���%e-�2�#}i���@B�^5�уj��\|u=ε���swf��(15��*�ڑ��Y���t�?顈��T��;ru4
�1�jػ�*?��@l��قH�1��󞾤�4��Z1<��?�B��.��jO�����)�ټd6�����t:m9���窍��F#f���,��w44�).7��#C>ʰy��##f�}�|L^�	V�
k���l+��%L�Ӷ���6ښuz�����ue���c %���)���0Ѧ<��x<5�!�f���c�������1Xê	��SV�4�4Բ��^{�O>���914D_�:6%��雉&��%ǯ�>�=��jQ�l��M$�����	��ǜ��p��=B�GI(�KV��*z���ǆ�ɩc��9�o��ݞ������֌����|yD�=�EL��Z'i:a�1M}KJ�?��H!׵}kl8����믻{��?d��i��{�/��C������F0֦j�����?�\�7i������5��	��Mcc���"y�H����PcA-!�{	�8�h�o�;;;�y�MN�/P2l>C�P�3�Ծ!4��b�`3�CV�)}d�'�4H��g�5�~i�1(���uZ�����>���7o�d2���j��0d�ш�(zps���(�F�J0IM!D�Q�씦ID�M�5���G��2�u�?�����-��:��o�=�I��K���ؤhQ��Ib��d�����K��%�u��Δ�*�Ϝ�]��#�9's��hރ8��
w���/>g>����a}|pz�G�9�[��B7�>���6i�fd�D�֭���K��9��6�"G5p��>����q1?f�8�i�w	P�b4X��Np��&x�:�Q��ط^g2������[�n����P-*�T�<K����a���tJ����k�k�6�k�ܣL�?Jm2|}Y��t���\��n���b���b�QT�d��z��������Y���{.�Ϙ�X��Q��s�w�i����T���*�4̐'���IڢVf��,�yU�3��u��9jr��r�����NL�80XG�ΐ��)RhI|^!HlSI!�F/��81}��;�.R8�MSr��^�Zˢ��b������7�`�X "�f��-��� �U���	wՈJ:m������A9�8g:��'��{����o~��X!�)��lE���z?���ͳt��H��g���MU'<��� �R�Mc�0M�}�6�Ir�:���rvv�x<f{k�FW��h+�8$��U��ǧ�/`<j鷼 �x��7h��DD�N�\�牠�T�Vz��*�:ùTT2������cDb�:���"����(eKW�qqq�h4b<��s��/EQ��̤ȹ�W4ՂW�~��C�����;�Ai��!���,F2��P��d9�h�+r����Oy�w����.�~��i�}��%3"��7��r� /2�s,�K��a2�є��o���8
/�P`���6�tL����<?/j/�\=�X�HUG����Yx�'�ߣJC�RH���M%Հ���!PU�шpnd.;5�90�F��;;�Z/.�*0~m��;��FM�S��1C���Q�*X�#M���d
��H(PM)L�9j"Zg�=֮1�A�s��Ⱦ;7UE}"��1@�$ǃ%D�
>�I�+O+ד�c ���4�Q�B�TƩj�e`2�$�SV&-Tc�em$%�������jj�1�&�z�'�|�/������є/;��4��}�l0}�u�M)6��o �������38=9O�![�rA"�jA^��.�����K���xe'��+�<�W����yxxLY�lo�r2��d��*l��A���/�ě�9S��bLd4cd>?#F�2��������4$gOk�@'�mLj��BĎ"�+AXGT%�@f�I�8=�9��t�<Z�8���ON��~��Dt��d��vm_�]�ܽ���ng���
���!�jko���bqq���HY���
92"��Ĉ+�;W~1s.o#Sk��r��}�D�w���b�QgBPT=���Gf���.� ��D�uf�1��)��TbhpbPIE ��!�>`2�8/��i�e��%��;�� �Tu@LҀ�@M�l�bO�>�+Fi�M�eY�R��c���8�O?������K/���8��g�/{��ED���{��#�n2�F����9��޽����z;�!yF5_B,g	U[l�f�����_����ې�T�"�	��TeHT%���t6�Xt����o*���y/׷=!�L���,K���HӔ�u�d��e���5����]mhؘ�����i�4��jA�@̦����]f-��kV��#՞�vm/�׷]U�1\�e�p;ϳ͞@�Y�X��1�A�TU}����ON��?{f�/�(6�m�bl#"�����L381D�k��✏>|���}k_.�W+��QbML��;�o�R�C̞�Da���e]�Tu/�m3�3��&���j��0T�Gu]3�����{���9���a��������g6���#b���]�}����\RUu]����O���S �˫�rw��� �qA�\�4�@�T,.��O�WDٮrD�d���>�z/�ʲl�w-���ޝq4>0�888�9��E*�0�~�~�!����[=�v}K��H����ΰZ����g���G��%w�~Ip��k��9::i��5M��*�
`�!�P.�|�f���<MN����d�x<���L�I]c��c$gwwc`U^�喦IrV1�)�l�Ř��X�\�ָ�F�awk�r� ����M���9a���).˒�bѷW792�	�k{{\�4�޽��⣿zO�>����yHS�g0VԊ1��)��{��w����z�c���=��W�FFmQ\�DH���N[�,I���L�,��pbhV�|�q���C>��"7�/K���'ڔ�M�����(�jY��S#X$Eq�U]᫚&�ӗK�UU���!�oW&�e�{��a4����*w��q�rY����o��EU���X$|�J�z��p���e�"�-ւ(�� !��^7�>ǫk�?�u�W�Ɠe������ۯR�%���#��Ƭ�ˏ��w�e~r��"bD��Lr�o�U��y�l��Eç��\R�O(�r~|ȯ�����X2�pn�b�"G��ܥs���4	g��"�o�m�c�t�у�Dk��L�,U]�\�S�Y�D�Xk�&G5j��E#B���qD�4U���A#�g��k)�N��f�v����k�8��ʲ�����qxm��U�c_�{gO�?o����~�b0F�5��&���n޼��ō�)ҟ�=��w�������)�-�<ʺl��1�5�%���5�bI��3?t<�x�o�ۭ"6��ǋG�9,��W���8ɋ�X��M]VU�Dz��\8�E�C�V+���\<M㙟�T��P55�npy�"�F�bZL`*� z�K��*��>Pi�f�RU�,�X��e�ȋ0��y,��Y�q)�g���dY�V�n��B�W�$����6�Ʉ���s��O9?����b�%��CįR��u�Z��zYQ5�De�8C%#����/>~���C��h��̦	b@µE-�l����}� ���Quiq�7�|�;�����cV�c���L��V%e�b<)���Q�d2�ڌ�+U��TR�dY�u�H$���
2��Z�=�1_��>p��.?��_��_������Š�9L�1�u�x5��ڮ�쉩�+
q������:&�K�cH�"W�5���S��oϞ�X��k��Z� �HTU���|�ѝL=b��G������:$3HV��Ħ�g0i��M�n��ih�y��o���%b��X���w sC���W`\DB�$s��ƈ� ���Ȃ4�4�@R�h5�h CTPb*&�*�T�8 �4uE��T�+`MFf�����p�����E#6kٸ��9HQ�<Ot:�ł�GGܿ���!�Zsc�(�E4]G�,����t9��H�o"M���fd.c����(9;:dw��l�x��t:�Ν׸��Ërp�6qB�b�6#����c���x�s�h�Ay��7�ۿ��|��'���s��U���kϲ\`,WgL�c�[3D�ղ�,=1���8'+F[$�-�Q^P�9���9��;����bvp��;�����Ǘ_|�~�#�#�f�Nߵ��ܷu�$L��w���'ڷ�1K�y#��c��2��o�[�N�ט�?{f��v�:�b���*�X��7:��|Sш¦�}І�dy�Ү��Z��XMU�Q#<j�t)�0Kǟe�d:����m��2w�0߾j[�+-�#�Z+�#��k��P<!`l�o�<y�J��u���I)
�!�DJ�V5�¤pX��@]�I�t�\���U�ˮ|�Ҹ]�9�}�z���)���dY���>�W4�N��P����9�t�Sa+w�Y>�19���h��d�l6�ƍ�e���)[�F������wU%�e����.Oc�Bh��=Ս1���͛7����;�&PW��Δ�����7g<.�
G��M)�-��	�%�fx��N��bB�;l+?hPʺag�s�/jƣ���h��rō��kQ�k�f쫜��c_Okݤ�Z����c�ƈ���Bhv�>���GnϮ��\�&�Fk��Թli�� ��4*D�Z��0��n
n�U��S 27�p��h9PhkNr�VI��AD%(fc�G{,�����X�i�@;�]a����nL��v��k�1�y5o�,����t��
:'�;��HL�A#�2�A".��?��Zub]�2�D��q3�����	�⮃��n;��x]{w�Q�z d�fL�H0�&V�|L'�r��9��.+�嗼�ڏ���f[�ᢺ��k�1�@�R��&E�@�b��''�l���MB��������bl8�4~������t:��{wy��O�h*��7�M�Z�@�'9����>� d�\��_-ɳ1�2�8�|�v~l��y�f#���!8�h*"ڻ���N"���=`���c2��뺯�"�7����2��Z|��0����ވ�Ez��L�#���YY�U8kɍ�=���>��|�/��ⵢ��:,[z�W��1�JQ3������ʠ�x4cȓhyb.,�^�~{�=ɋn�	��(O�����/ُ# �t����ߴO�� R�} 3Bp���E`���Q��&XS�e��UxW����?�y�{��5��OĞ���{S䙫�1*>Zc��[b#q-���UX�a�eh�^v������.��[*i�H���ገQ0���V�&��ld�1;Ƣ^9�H��!�n;,���E����988`6�Q�k��,���L��~�mn޼�;�ï�ׯ���ҴE�`ggg�6�,�ma�e4�A"�/IIB1��\I<b4U���k�:M�}�1B�5>4L�#|�F��������`2���$��U��Q�o,1
D�c�T�h�(��`\�ƫFa2%�ؤIAfZ̆���hDY�,�ˁ��z���i��4Mr>��#�Yv������o2��uXG9�e9�*B����},Յp���gv��E���K2.�2hC ?j	��ݴaz���u��/�Jr��].�����I�52t\$����!JE�%�����?g�H���h���Ísꎣi�6ř����-N�N��S7%M�B`kkь�?��w�}����_n�\��'PV�1�,3��cb�+���Bւ���K��ڳ�͋("�!�,��|�޻�f3�g�̶o0��߿��=��%U��E�t��6�x����o/��yJKR뀸Q�~z��,k�j���Q�1��.)˚����_��8=;&9Ǯ'��a���x��]!O*���Zi���x�i �<C�Xk]�qbȂr�!F~�_�������OĞ��3��7�I"�1���E�T��=�${����m�B�N�l�L�pi/n���f}�YqI���rT"Q"Q�zNY/�}�ƒ��SV��ƹ���h��|� �EU�V�jA�G�N�Y.�NJ�+֦������"b�1pcg�<��f�X���i<(�3v�ʀ�a4v���INP�K|(���
Vobrh�}/��M���O@TT�s_���rt|�'}���vw�x��g��z$ɲ;��9�^[|��-2kk6YlvOw�C�%B"��a ��[�#�A����y P�<$j��iABJ�fi�Iq��j��fuwUu-��ofv�=Gf����UDdFd�/��%=�����=�,���ob����loo��u��޽��l����x�Z�qU�ށ\��h�����֢1fޖ��*E�r���>{��t�<O��!�������-�d]:��xɕ�=ǵN"�u�:bb��u<�����t��2�܎Sd��I �@4��j�U=��dǵg�*��tQ�Fg��f�?�"@Ϟ=�t6�phaB>L�� ���SXAVa���H]U� �AQL��_$�'*��s1���Q�ʢ�?Z� I-zY��J�O�0@N�1B�D�"v�	���w�q����CiP-k� h�	�z�]0��5��@9�FS(����� "`w�)>��
U��ܹ���h4�[�-�R�4�p8��=�y���~}~��ԲIm;�v��j���i�����柟eOD�    IDATB���rV���^
k�n����BT�bTUk�s�5�P
���lx��A���Y������ z  2��Pa,�)�O��	x$����&��d콟W#��*w�2����X�9P�
Fl��	9!����e	@��C�Z�n�����F;�L�_�V����PI��=,�1�e)����
�H8���3T3f��k*(��H���D���~��;����7�	�����!�=|���;��U�髯��誥����4 M�
�bŬB�B1��5��0������a�;��$�F�3uol� !�ab	A�6�k�I�=��pi��u��Z�� e$V�������1�.��s�6��x��9��)� ��|�s���e�䝄��'Q
@��a��"�"�,S��͛W��v���W�z/!8%�* D���(����m��������
ۖ�*�8Lq��w���һqR#Ԇ>�b�<ϑe(|T�߸��~�����;��t4; ��\=<�H���$I��iӓ�����|.�=�L��o�7n��H����^�\�=�=���;�ֻ����|@ݲ�52$��X�D�u�PS�x�������b�B|�?�s����B����y�$"F�H���3(	�� �`!^�� �����E�S���ܓjc��U����	Q��!��7� �Z���Q�T�^�7n��t:�{�F��"��hpG�kD+aԎqQ���2�<��n���d���~`�k�錾�z�*U��V�B�D�(s��{�XΫ[�������úz��W�p+颵D��AF��`r�JE�;�o�w����.b9Äj#�(j� I�y�d�=vvv�OZ��s�!�j	�,���E== �L&��X[[C�� �3��>���.{I�!1)����d
�dpFPU� ��B����AljA�3���*�:��	����g���� ��>G����p�]�k�
H��
��U���A~��c ���4��i{~�6��Dh�Pfn:�� � iB���I[lT5������1F|��g��f�y�fc����u��\�H�q�ڕ�"9Q�(��T�bϕ�1��_��\9���'�1�5�� �����g�U�HI�`�=�u�I3�:|���"�<:�+�$I%Yr���4�줉ʫ
-΃�>ŋ��X��D �ß�uv�"���XW�Ɗp�7���W��7�o�c�����7Z�+�v���4=�Z��m�/�~��q�1l�s�w}�[JD��p�U�M���d2�͛�P`2.����|���
����A�A]#r�Ź�q���n��|���`!�����)�ky�Eч6�#Me1ڟtt!w� � �}����X��펡	o��%�(s�&4���RK�4�i�@u��$I���������N��أy��a���뻼�Yu}~.ڨ���q��w�ߟ5�q�y��H<��,?�X�Ԍ��M V�9��9�z=$���g���!�4�T�4}eP\]���������������w��>@������.�{�ۿO��v��kU���p,�u$t]����q��[���)qD����S3�xv0b�x|S��vt�\�
!>/.�-b��x���,��v�B��ԤU�DX��a�����h�V���b|_Ǹ����o��Eh`�~�Wu��A��w�Qp�kG,���i,����݊Dn������PE28*A����=�TM;2s���|Z�r�Q����K
��*n�婳[e4.m�1�)���&|׺H�̊[[�uo��s,���풂��L���cgf�S��f�Zs���O?@٦��n�´��@���wtA�3?����i0�3�f1��)�L����N�
��x.61�� �C��$�a�۽`�K�Y!����D�Y��8�p�Ԫ�@�>t��Պ4��Zԅ��5�.Q�������;�����q�V⊄��ەK��g�R�4��o~� mf�ciߗ�3��`8�������sW����g�$�~y.$�Dishq#�ڻZz�P6����?��iM^'��>U�)�������VK�>����Ͼs�G銼�d�+y���n|J�k���|<fn% �"������ ��
�K|���WB�q(����"Y��e-�hM��Sm5w��@1w�&���%�>�q(N�_,�ڗs���^m�_�1d��F�Y� hjd̞E6F�����E�<�K���R�İT����eK?�t�*�r���)��w�X�m�&B�d�5#2}����ü/�m�ZZ)�>���35�_�֮�9����Oj�2'K�Y1	ͨ���Y����c����u����U۽�jl��܁��|'\C�UDJ���DpD(b�/���[�����q ~�HJ�_�I�6H&jjf�p�dBI-S�q��*�l�H8�����ڍL��H#p���o�OX^M�x��4V4�_'*tvWI�"�Y-hXT��"���?�&�]w�ͿMb���չ�+�C� � ���۝&�m62Q��wd|g�����Z�jL��͛�$�q���J9�eV�����d��{*a�bЁ�O�e����l�2{�bu��2�P;�z�݌a����ݿ���q�m�SH��� �n�C[���f�F�Jg���h4���*�𱱣�Ш�H��	��U�;A�0�c��W�B�������MqX�մ��!���D?*m�0�`�`YMa$E��g=� ���9:���W-�%��%�����1����6�+��L�W�%jf/Vu�0�u���s*��
��
�w5�F���v�e=����{Y�수��,�5*a_�j����*�j*lU[��P+,س鴪�9��y�?^��p�Z��>f �E\�r�"��Xq(�Z�k��}e>��Bɮ�V:�k���T�"E���8M%�M:E�i�􅲯B�ǰ�*=�Z��O���Hl8"��� \V��:%.y�����t�Z��_�g���V>/��W'��9�C�����Sc:�.��O�_��������ާ�9�ִO�_ZiѸ�	!ı�h��_��\�?���Y��I��W��G��}�e�h���[�������b�lQ��o����R&���E���Y��u��;�#/F4O&�7J|LݽD�:��\U3*]f����0�*�W���P��*���}��{ c�X%|��P n��1T�W����k{��֓��|�?*�{�Z[lO��k{�׿1�g�%��
�+Z�_,�Ԥ�Z� ���^I)k��g��(y:kƭ�N�ؠ�O]�j��j��HK�GөzGǗ�������B�X90����܁w���`{i&a,+;f>j�h����d'��%W�Qk��9�L�W�' Ai�gq�F� ͧ%�����f�u�o9.��)A�ny�_��<l��w(Y��4}A�^���h��ύ�6�"��`.��~یl�Kk�D:ퟤ���5q��l�e�:pF�� i;.�A��/�3�SEu�*5�^���5cC��~dO�^��S��#����֒$"�*�qP�7�o������yW���WM?��o�rMcu>�tJ��.-����x>dp��|���?�Ό�z�fَ��9p�+�̓��DPή=mO�����\�7	�FF��M�Ց�Tf{��RKE��:Z����<{k�����o�{{�B{.���vߞqU	�in�P190!΢miL-�O9j�a7h����1�}��z&L1�IF�)V�#�)����!��4v�Y�Wn�P#��P���%���.(���VCϕ�J6�=�T�%d�*�+�f����e�=k��Kj��צ.�92�6����
���a9�d����Cz2.�@^�QoP����)P�<+'��xE�'��=Md�;.K�E���x���l�HEt��p�!��O34"�:΀7M�sqlD������y���d�XN+�I��%�u�<�qve$q�RRi�/��4�ģ�o��XkF	�E56R`Vh�+d�K�-�t�s�S�6���mK������jE<r˳���C�,���\��P�Ilf�;�. ��g�zo,�eTE3"7��Q�Zьm��n�����P!P���a׶��G��3�B&��rK\������}�������GF#�����{\��V�D�Zp�/+m_E�[X���Xִd>��,��8呹	��l�K95�~���ңV��sqC-�H��fh�~����C��r-�����̕H.js6��S>[;��"�(hmB��%<�M��u���+D>����
�=�Ѐ�˱���,�����0� �o��D�	X���}+�$IIIk8�SW>0{X�%����_���˷M[ �}��S9�&S�I�������9�����sN���|��*!�4b�a���L=_9^��$��ys��q��b/( ^�և�>��d;�����d�E�T{V��Q=�r:��l"�Ft[Ă������9��Tg��/�����'����!�Yt����!�YMG2����p�´[���QDJ�AM|J^�1o�}�ƃ| 1'�!�7��G�7|/�X�C$L/��j?F~��ώ�'�IY�gã�R�"�d�d�ꆠ�:Z�ĝL��?�}zS�ëq� X���λ�VZ>-�g��Op}�S<��	Ƚ��611�LB-�K��v7}��탿��1�qq#�۝��]��*y�rF1Dg̽%�ʲ|�Tj�@����z�\
�~z��66$@Ʊ�DՒG�_(SB�d\�`2c�.0�=|f߳����W�^�j��[L��#g�"���t+�X0���˚� A��3u��L���|�j����C!�&�t�D>,�Z�t�������)��I=��C@��ǥ;��5�}:�}�[�h��B�.2�.�AR�y�!n�.��.\�X!=g2�8+�ThO�Rj�:�¢1k(0<���B���E�H��2�!-%BχŀZ�S�h�W�>�Y9��_���$�i��o,�=L�y�Il� m��8d=F@'�|HR�`	9��P��{��8�srѥd��t���\�ċ�� ~X��ݝ�3˔0�-�͘/�J��O����x��ƴ]��[_��G���v�t!lUP�I�2�u�/D Ք���L��(E�LG�7����bZ�\���ȴW5�,�\[pر����qد.���y��O���f?l�o=�~E���}�F�����>)�uS�e�>�����sڨ:TH�_��m����E�$:i�]~Ft�zҸ��p6a�I���Z���:u_��,����h	�A~sbR�U���~9o��E�uN�g�������&��d$R�4E+�9R���Xȇ$�/��W[�^wMY ���DY��aG�}~�����}̓�>Қ��o�tn��'6�.��`q@��4�@t����<��J�f�rMو�����1 e����Y|���z��{7�옾�Z�o�����:G~jK�6����TM���f������f�LF@�D&lX�j�1�3��Q��NJc��+1
�EL(�Xj�4���_l��C2H�-v.�������x(6���N� CJ� �\0�Y~j*����v��`�n�����3NRlWR-����������T������Ժ���WeP�DH����$۵��K7]�h���9�5۠�܊�����i��[/��.?�S�0���j�~a�FY�	<�Y�kGƠ�?��+5��@|��`�ge��`,VN9�3���$O����_�����q�Q��0I��Y�_&R'��K�>zF�
Y�T��i`G=�ĥ\�`����~�x�Yd��i]e��� vB*5�$;ﻩ����\��$\a\�� ��4g�Rj�V��\#�%%�@��|�P#)��q������8�W-����q�p$,�"����%�$�/�#w�Q�!���>���G���ĕ�C�~��'� ��޴#�&p� �zg���S#\e���!
��s:۱Hi���DT2R�������0��1���0d���ԋ5|e�2tvn����������������d����L��Z��2��1nf��CK�hp�f	;$�K��^�W�9VQ�1��r�u3�u�;��S��(&��	je��A��/_��Ӗ�Ц;�eP��U�[��b�A�d���1�����5	<��g-ԕ ����_�x�&���&hu�чe��]Ģ�?즽w��:�����]!� ��7�֎g��wGPe�M�����8��׬>��f�P��G��(����Z��k0�_��Lw�����'��w������ܸ
�gh��sUceLM�f�M�5G�g��ݙ3=�!���Rm��v�K�׿V���%~0�VPQ������P1��f^�,��� $hf����,{MkۂA�?B�y�X5�9׆�T^��}���SAy!c��Ie�������,��K'�6LY��2�z�+��Eمϟ��Ѿ��<	Q�����A8�1'�+��j{h������2��K���C_�(:o����������=,~���X�o�/i��~��ۧ��sW�a�`�@��M�qF�u'+)郎J��	��n�;l�Q������7��P{�:�H�-�Le�]���?����zo���@#����x����X���GM�4+����99��PX3O]���P|�Z
V&�n�e��Hӵ������.�ҡ�`E0+�i��0�}hq�.�
������0�L���n���/󾦫Kv��]��;���c���ZON����ޘ�������)�Sa�S������O��8s����_��/��������D&��v�[��v��{���|e!HN�vWx��3�P�lwq}�v5��V�N���-�T1����7�w���SߚF��{[%�̰x'B,^�G���N��UZ �����A��q���^��
�)�Y�6���Ͻ� [�������zݰ��	t0�QP$�W�l�lu�W������f(�)�Oo,>E�!I�����!��g�bH=2+ǚ׳�Jg���sC�e��0�)G��2����� ��6K�ڭ�P��;���@�2��%���p���~9��?tn7�Z����m4q��ˇi�\F���PzׯT|�\�J����K ���p^�H��͕����t��Yā>�qk��d�K��&SX���Я5����
��x>ێN���3�!
�Iy��oA�M>A!���:_L�w��}��8���H'�
r��=T��U��B9#)o���:��'>�;�)������z��Ҥ��!ɆA;K�WT~V� �VӀ��u奔T�[PwY\���ڏ73���A8,������i�!>?��r����n��g��̼Y�� ���qbuZ%���4�){�?T�@gQ�4|¿ո��`���c[V��4���i�s�������o��/�,�WN3��C���F8#(�l)�*��U��_u�5nZ��o�c�Du�&�[�z��O�/���}ă�ݏ�}y�>�?����u.ՕR,�1���N��Mν� .n�SqG���d�(�M�$����#^���<<A���͇��n��M������$�����x),����"L$�V�g���&�Uj�؋@N�U����������܌H�s�/����\�E�����moΞ�˓��:xm�WG�83���Y|�H����;M�:JU��r3Ҙ&�@$��Ÿ�y�a����2�:�4����%Ȓ-� ����tb�00��
�+��!�ib@���{i����ܬ�,H͇�j;XM���I5�?����@�tq0�U��Nx��i䕿g;'f������;�&/�֫Yx��DG5�t�I�p�;������e��"l�}�]�b|[O*|2��&׬Xo�"d�H-�����o[\YBv�|�o�7,�(�sh#2�T~�ڎ���3Ko��,�IH	cr�C=\n̩h4����Dگ�x�����-�'�"���k_�ٽ���"S�k�zW�6��ab۵����fK.�I-o���X7�)ŷ����U�-��Z>�v�|M7Fh(�U��tj\ﳒA!be�APt{�/~x��Av���=�^�X���XL,DG�'���G6�8q-�̧����@�m�0y�^K��������EG�uM�~����w�3a%�������ƛ������LO�g��n���n@*'�Sv�V�I8�]���.&NǞ���ã"��/��ؐQ$$k��s���c/���(x��J�յ�Ⱋz3l�G�RO�j�Wb�(�#��X���%A����o�&��s�b�>Z/�.�h�_��W�g�Gy哒!a0�R����7�g ���� �0�@�,�n�"tg���������)�+��5r<T#��ߔXɵ)0?Bo�F^�-�`0<�@�a1b���ƣ���i�D�#>g�1-�膷��j���.$�-4�����}�Á��{��Y��N���[kC9�퓓�	gj��FZztZ쌼���2����G��̗���\l_ϣ�߷��'d���Dh��m��0M��T}�5�#J*i�J�w��Yp�%����k�5��9^\�O��U�rt����rKK޹�Pm���&<�(v��+t�2<cJ�Oƴ}���9fg������4��j���ʚu$nG�
��џ�O���u�aJ��
��v+�O�GQ�����TVU-H��)d��֤��*�n���̳k�*�T�Z���.�5�x#E�4�c���L���I�|�*�/[H���C��G���^�*H�'ͻ���U�)LC��iz�q1C��o=�e�o�}2y|�3=�M��U�QT�����ݲ�L7��\M=�zmXw�c�I;Vj�P^4��e�3�S��/�Ic��`:���_���h�~sq������u�ϲ3/����v�<�?�NED�+?Zߌ�s �N+D�I��(�wPD��-+�$|	Y�g�$6+��.?�Z����t�3`��<h�Fru�E�K�qÚK{w鞭v��
xF�v	���"���P�D��pJ�Е鉜i�r��g��&��Ʌ������pe����'�w1�A�X�JAV8 ��4̬�����O5��_�89�?P���w�c(��f*�3��^I^���L�{M���
ΜO����n��oϪ�c��^��Om�?[we�v�6�������3r�w�\���l�}F����z��׿��_6,�����oq��-N�O��	���&j�S�\�Q��N[��X�j�xवc�<|���UИg���]=Y�s��`Bx�56���l;n��κ\�9��d}�/�'8 z��MNO����k���$B��u�qiC@��%����1)�F�~M���A�����@�����`z_Cn;]�wI·��?I�`\7�������E����d��gK�����1;TnG��r<���J���H��Ժ���y׽��j{�H��(Cfd���o�K���;^��9M�@�CS�����>�~n�q�����S蔒2&V���1���^�e�H׍rĵ`^����M��1�������z��E@Δ�-/0c��d�P�7EM�����w\\�h���&�����g�@{�ȧ�5�}����:��4��Sf����f�.�+�(�X~�/	��_�Ǆ��lJ'Q�4��18±<��+�_���	��<H���qo#����?MŃ۟!��7G�ɟn����ݽu��	"��m�cO���[�!/|�����6�;�
������y-��T�v���z7�ĳ�;��G��CPx(`�*!��yY~e>B��	��l�����{�H�@Ҽm���r�'n>�;nő����0"�F,��@��򗑨�Xh����Q�T�kZ�f�Q�Ol�����I@ȃھ���$�{� Ʒb�n�M;;��@���xOk�3����z ��o:��u�a�O��1��d�1gk��v�J���|���2�  hen��86�sJ}"\[.�+sL���}]�T���$J�+�3\:S����{�*�	z"�8�|fA�2K��.��긶����ո�3�M��5�e�x�|OƝ$K9Q���.J���F�6��6®0�>�
�؏ �{Q����q�oh���!M��2�'y��t ��V���Zy������򢍛����Vv��L�� �{.�3�7��� g�1y|��|g+W
7��	���xh*�s��0���T�w}� (rm��ӏ�b��")��k����JT��p	�H�����8 S�9Z'��B� �j>�DCN��J�#Lp�HlS�$*�D�'i�� ���#q	�$��W��G�ogfE��w�t=���yI���dbb�DS�c��9g�˰��n9޷c%����fb�(�w��\9����n؛��s��zF(LV�.}r���^��^�n{��vݴTX��jB��P�gee�e�@My�m;�ω���)��xy %�������)}�JO��?e�`ᡰz�,�D�VZU���o�Nd~e7��F�V��	�./j��ܲw�W�դ�����񅄈k|�*bb�+\T?�˟@E)�\y��h1�EB��'ؾ|Y{ۓ A���Ɠ���wϽ2�F{����aƶ��iɘtm�E���s_�&�_�A5/[������o�h��hp��ϹJ\S���7�";���ʡ�ӝL����ʙT�����L6R�I��r���l�?bA[̘gY�
Y�7@=s�P��Dl��ׇZ��W���K��!�=2�&1��G��6����h(�?��\�c+��R*9��)#�H YU��y���>��E_;���  ��f�j�e���Yョ�ޡt�x�_=|�r�b�
�7���T|'����G�
8�E�,^-��\����
.n�ӷ�5�A���z_!zSO�宩�f�I'":��������H*S� 0E���?�}��E��_?�U���7�W/�Vqf,b��L�4є`	M"�/,|n��	�/**��f�ṷ}w=��,�+fS����ᗛ���K1��"B	�ݎ��5Yw0��L'����:���k���`ᯮ6�4�W�s��X^��Nط�ѥ�^T��vPSp�<� ��iU%�����g�MFu��4��]cg�-���iZ`�K�B8h��`�����u�&CJ��a�q���x���b�q�$�F��]QE���F�A��T�́��2��F��F{��i��l���/}�H�&x�@+0i���s5(�us2?3r��@F�B(G�o�=Ώ��E*��'���Q��SǷ	�����Z(�X#�"6����y����S�IE~J*ݤk�O�t&0w.��O���(ͱ��0��6W.�A>�����J&��lM�6[v\\_{up��F&�A��@��ꭞ�,#�M�� �W���e������c���Ǥ���3�H��j��Bz���NҬ��v߾g?�:�N�l�W�U.���jp�59���
QMѶ��*�%��x�cn�u���"j�<L���гhtY�w*��$*�B�Ԑ�RiԬ�(x���hh(���vu��͏���rۀ�|��_���%�<V�JI�L��7_|O6s����mЗ��;1L���������㿖�{t�>�,5��?D	�{��Y�E����RM��� 5 ��܍�E&��M���UC�!j���d_z�_����ƣ��`d/�\ݭ�_7�v�q*���Yt��C=ӌ~w<Ɵa٣5��5!3�Dj�A�J⧃͢�5��8ס���yՓ�X�$$Tl��#"��r
�?v��5=�c��0� 0��!�"�ՖI���í��)FS�&#��CC���YR�r��-������H�\!�r�9�+|W;���h�2�j�^���ү�̨55S3��x2!�y>f�B�~�@�A2�,���0"�h��	�����IB��@Q�v]�rGH5��eZ٤�5�����\�����E[���2�j�|�A�k�R˰k��0u�3�A*�r��}����+�߁���3m�-���_�OW6t�����7lR\6�gw
b�q2�tJn�]*�X�G��;��=<R��~:;s��q��D@�8h_��10��1��y�Vl��.Q^ۖ/���uo��s��מ��T	��xV53c��)x�e�W�V��A�� �j;�[�h�7�(xo����5LEVk;��u�}�����<���HI�
�Ї�^�@xq�C��d��8/K��*q��=L�pkqk��g��g�Bo�C�k�B���Y���G�����/3D�\��v��}�cTs�"�my52�M�@�T����Ǽ�܁-�ʋdݐ����=2��v	?x��g%�ӯ�_�\�5��#��gU�j)�ȋA(�yS�g�l* !_�]H� �i��S�qs�,��Od������e-�;cFY����'�2�j�޾w�x���7��\騿��ԁ���V?�.n\�s�Z	MJ������5�I����>8��B���w����7��IOg�O�pG+���A��J�U�I����`*!��'�G��Y�p�0[�[G�*˅�}������4���1���N{����
_�Q�q�`�V����"U`*��g���wm�����o<�nٱ/in�&{���_P���&�Ʈ��P"��bg��(xڔ�B\FU�s�m~�����n���I�'��n��|��#U�<�>��T�-K�3��Д������SB
��<����2-����Z.���0cY�hZ��7�m[���X�K����͐�iu��铍$~Ԥ�Q���衆�M�S	(Dܾ^޶6�0U�^%�����'���n�=�0=N�l��T��\L���$l�����bM^<��ʥ_�#@!��&�(���8[�ވ;��PV:�1}�Ye"��K.�Sx�8=��
�<��tC���4��İ�j�$�B�|��	}u,A�����O��mc�B�T]��;s��$8(e��Z��j?d�q��6ӌp�#��\1?`l�^#��yÅd��Q�ح��Q��R)�g<M�@�ϵ(y�����s7�N&�q-jY�~e*�,@!
�*"$�I!�/�z5D9���f�ņ�l�Ww���68jڝ��0�K����*�Y5�O㨕*{�� -<�&��dX�^fs�:�Q�����_��&Fe�fğ�J��ۺ�I+�rp�^�܉�s=e;G�����`.�
w����J��q͵:t,l�P9�>-ڄ��	����7y�o"L�j[:���ow�s�\������HR����K�#&�K`N![^�C��LȘ��,؀v�%2$7>U5�������d��gP����Uu�6aF��J^� u18�����^�uTDxX�b�/�U}y(� ��uh�.��if��J��1P�T	��CG�ۤ�����*���M�%�Df10��E�����l��d#���5�������
c{�<5zW	����Z۝�iB�#�X�H���	--���|�����a���0o{�$SYm�kk��Jo�%�����
��Ad1�d'�{ƿ��g�L�����}�@���	 ����P\��pȎ�k�Nmuz�|��N���wnd�l�5��-���D0�%�L �T$�J
1F�%�����&���mGx �ƚ�հ*TJ��a��%?��SW	��檜�Y���3�!=�^�_����9�Ʀ�R/ɊO�vU�v��Y���K�߰Ʊ����E?iW����֠�%S�%P��Qa2����#a���#��uA����_���[�{{�Y���I�Gc�0p��۵�KX�嘼1�j����M�n��rYrl�����C�� iZ�*�o"��s3Ɯ����C]�������Y.�����=~��������h��h}���P���r���&>B���D�A�?ov=� &r
�o�!=(s|�g���,���ɀ)��A�jր���xr�Kޗr�!����~�u2�-˘�����y��g��66S�>jq���SaIY� (��:%m۪ʔJR�G9�X$b�ԩ~�K�Z`���[*<���W�D�-j
���^vĆ�!��>o�Jph�Ḛ`@��,H}��@�?��9E@'����g�+���HMU�.�)�5c����hC�<:ں�b߽i"��q��3\�h�����{��Ǖ���#�� \�~ؐ��U���zv�V��~�A�{�_w��NrM��&C~gn�C+Q���b�)[1�HD�G�G�΂���0���c{[ۢ��m�X��Ȏ҅��bP �Hi�Sy
�;9��"�W~�	S�
���m������A+j����sL��}\��D������{k5 yxx�&�?��o0���ݧsl�X��
���&Ao� �Y����7���:���,��M:*���פ�Gs��GA~f�Fm�1^'�42��yq����d��Θ k����5������[��,資�&FfZ[�=]Y�X�*�=#�r]�5pM����-�y�嘟�������w[���ލ?Å�I�>��(�hJi���3�+EjU�ɨ���'J��%uѦ��Z空�����n���eu/-{�դ#�5q���7��w�/,.fD3�`P(E@�����ݽ���3��_מ��k?;1���VW�2�ĕI~�p�2EAO�~2	od�?���'��N�+��܆r2�48 �~� A�%H��1��1�L��T�֗a4q��~�r�v|�o��4!T�tU��GP˛1_�؞ߞ�w3U���ԣ穀<Ec�"��/	���P���al�T4E�����ݴ���ܘ�5�1Y��+!z�:���ɋ&:/42)�����V��3�t�Tj�*.O�F�\M��À��*���L��K�*�w&�	�[l��H�����7���W(�B��?ц����X�w+�y��#�)O���GQ�>MSCq|��GI����M���뭨;)Щc�E�	��j��[7�Vo����	��ʯ�{w���b�C,�l��E�����@�3��j�-X�~��_����!��r���3Wq:�wI��7���Ns�|I��^�}�dO����$8�r��v�̊�H���p�c��7��O�+,��Z�;����y�7LN$�K*��IHF5��|�@<?�O@�8��o�g��z f�6
�����'.���/S�Ô�l����<���;ã2����,£Eb1f�V`��T����7�)�7�2vL���+��ŏ �������xu��@���w.�`F��<�$�#�h�:U�&����M O��T�Ğ=#�̫H�LE1SI�k_���}>���H���=�g݇�u:�ɔ�
���}���,���w����B�ϻP�I�*d�y�\qX�^���to�q3�a��`{�%���z}���sWmt C4T�OT50=LR��-�\Ǐ����ͩG�?�#�J�ɦZ5A0�t��F������y4)`p��*Ԅ��{?]Yˬ���W���ge�T{�uv��g����t9����˄�5:�A�^�=�(t��beK�4�l����u�6�j�ءL@������eU*S���vX����d����OjS�S3�L�0�:O��"��=w/9���~6�CJ˭�Ic��o�`z��{ϡ�M���g�vE9���wX�1�M�!̮Pm^ٞ����L&��"c�"�t]B�j%{h�����Y"qlG�@"���o���e�Q�b%!!!FM��D/�)�9���(=�/p���+ ���ږX 4`�?�����e�g�\�i��+S�k�u����;�`�.��Awl�D�`|L�Щ5�
طBƙ;G�׾g��G�c
x7?@.�Ն�~���h:����KjKYI�/	ɠ�H��H��S�҉��d��Mj��9��
��v�Cw�JQj��w-?�ne�=U�3T��nF�	>	���@q�M�b�*�_��<GlO��>����R��iQ�6���?�N�|_����9��顦 ����R�*(�f@���Qڿ��6�έpc��D�:L|�o�P�6�|�{-�y#;��Mi�3Noyx������k�8���$��ּꜯ�w���k���B	1�#Bm	��qp�t`�e�P1d��v�P��5��	�٧z��Y�)X*��bD�|5�����3��gS����j�Xb�z29���Z����"A�����7^!��M-J���1u���4q7����&&vo��W���~,&1߇ q�u�l���ۗ'-�]_�RF���Y����H������{	��3���]�yp��lk��g�3��$�[O���OJ�w���k��x&3��q�H�,At �`�a!Fb�[J���z��ũ	|:@4G��9�OR��0΀��Ҥe,&�8s��C��^��;��@ׇ�,���D��I��@=�Yo�q�۽��ΐ��`(�sG�{��նVϗhv#u��6�.�S����sU��^��X�}�!�I�O�Ԕb$� e��YKz?�̭E�c��?妥�E"6�� @��s��%=
����#p.�� �X��ئ��\P�aE �!����]���;�i5�m�e*�������Hi�P����b�3؟iV#�ts'��7�UظѮB6��lK�����y�M҉��j�Po�������������g�r:��f��8H�H�C)5]�����z\Cߦ��*/TvD�H�V	� ���&o�������?�Q$n�5�Q0��땢�
W�o�99�[7&��`������M_�
wy]#i��}2����v��PZ�b/^�ݙt�����yt�`$��*sS8���z|��I1Q2Z��Z�VG �y����vX,#R���fX �B�ŤX�X�?�	���x�:���N������p㕈HA	��iw�d��t�
���u����_�\4�������^�	?�
�M�e�~�₎�a�ο�	��r#���?��x���x{{k%����:WDi�\����_E���5S�U�YI���/��7�L?F�8x�7t��id�Kf��]X�{�W�|#�w��Տ���B�աINT��ֳ�}�22!�Lma���~x��7�]>O|.�S�`��7_�?�?�5�z523���7VG���]dޅg����$��c���5��p�Q� ����C�a��~�i%h"���u՘�-f�z}���i� �����N�;�z�r�Է�pD� t<�8���XI��:��)��P'�	
#��F��J.�<n�FO�LN��bݢL��A�̿ ����G�Z�,U�����	�G�w��$�"�EO�C7��{3@�ۄ=%y��&��lۗ*����؎�%��]S��+c`�N�hy/�Q�?���mCٗ�)�C�&q_{�����[l��з���J)�H�d�ym�ˊ�(�
��\�&����N�)p��z_��V��~r��	�}���b4x����'J��I)�)���O#��$�\��=�m�����������m޶2I|��eϸ����gmfo��=nt��Ob��8���9�7����B�P�E�O�o���ϲ�<�ʬxQ�����g����ދ��;�������BM�kG��6�ӛ.tY~��y��}z(W1��5L^[Ȓ.��]�K����u����=v�(��p��uͻ���P�t1�ZE�!������/Q�iR��L"AwGKwC�������^�����ۛPe���M��`#�H�fW�
i%�P�����@e���3�W��t<�c�ˠ�0++X�y�����6��!�Gw�|� �J��A$a���>�v��d� ��#,,JQp��^pW Ĭ�)�����POu�Q�(w�pbޮ�ПL&�Z�(�&�����x�I@�Q���/�#c2�r?+����%A�rF�R����w�?�Tg�r_�������{���=�_a�V��������o�`��~|���p�����0�CK
,�����훷?e�*�K�Xʝ��.��E��� B��
��|���fa��#M�y@0�	�K�Y���w A B?�T���v�F<�K�$6��=�@:@�	V��o%D�o|r�ѡC�e��vww1�E�iǓVj;<=���w<�` lQA4�i�� iR���2�kά�N�"ů	�ϧy�Q�')�]{��'r��{��/�o����8e}����,C��ׯ�}�x�ė^'�k ��O"s��Q!����?��p0�z�G̬�F�b�!��捛���(�}�Rĺ��E����>?��cb�xHP���4d1Z#Djӛ1�� ��� 
*d��i��h���ܖ��/Y��� Jd�Z�^�J_gy1�O�OC���75̌$�VO��tc]t{����1
�B �� �Nr������DS��|�9���ٰ*����/�����_��{�����R���ܛe������Je����anXB��V�L�.ݤ�}�k���/'�����"��&��K7�����^f���l�|RM/���>���d��;��t�kr"b�I����Ͻ��7����6��c�i��^��ۛ�9礎H �Ci��	���pN��+A�����o�e#+�z=(V �'�@!���H�5 Cf��
�DP�i����K�C�Z��i�_`��}�O;V�^�Β ^��|�p.@��Ĕ�<u���ܔXͲ^Rh���a�;�]"�)�*�7��?�I����[��9��~�s_:7����)�YGH`�� *]�w�p���?V�S����W���N)H�3I�TJ�g����>�v���x"��>u��g�(�>92Y��U���gG�Q�^.���P'����R�͓��0V�Ƙcjͽ�[�J��������8�<D<z�>|){�� �d�<�)q:<\<�`f���wr�@��QH��
|q�;�?��F>2sC�S�ӌ�A)���p/�[� J��×��>e��$��
1T���DT26:)4kd���V�@`o�W��2ɏ��k�Ի�V��W��g��P�������vP��4���f����C2 r/;?�hP��I����1Ed�[����={��IZxo�d2��Yi�t�w����;���GH����؟������"�{�h��*Vױ_�'+�W�ui-m-��b�r�#�p��<����&�1a��~~CSt�/���ʗ:%!"����D�Jڃ��o9sx7t�p4�s�C�Z��&�{�9�4i���q�� A< q�}�$ H�$9�Oi)5#�T��Q!��M+WlV���{�>��}��
�4*Y������ �2L}�x�2T*ػi�6�֥�W�+�[���p)B~2�j�?Q&aEdX�`�ɴ?����&��I����s��ō7�Ĵ+���y��\�?��m��3� �<����X����8{�,�y�\�y�|�<�r���w�܄1�Q�݈/����')�ە��+�< �k#8 ����Ȥ����СP�#�w/F �F�>��H_�^��\ 3��Q�0 �p��H�N���'ȳM�g:'��wΏ��=���Ɣ}3�� <�T�J��t���e@B�����Q�"�(HP�(S��?��2ڔ�ZUي�D�����Z0�MgG����V5+N��~��5vww!lmmaV��Y�&g�v.<���ڤ�6�z�hU� ������/��,��;��;�i�,�2%�u Gb�s6�<���!tu�g B�����D)�{�����Y���f�CT��t6���;�B �}�[�����5	}(���q��*O�.�N������Qณ���;<
����ó޷��]�J?h"{�`�Ƈo���so6����G���g�I��$q�ϒ�F'�}�[>���r���R��|�����}��خ3��ѼDf>-)?7�z����;�=��,Ͳ�F�C��J�� �B$"�
y�� � �uI����"D*(f��U@(��(&<	^i�"$��6+�B͊Ib�*#���H�Ib�!,���Դ* �\� �Z���Q��ڷ~���ج�1KD�̤�Zk=�I��,˰s�^���{�Lo�D����?�'��]���硲E���Rʧ�F��P���]���1�J A)�s�Cu�N��h��H�E�[աýx��?�XMY�:�P�^)�%L��"�A$�.H���A	)�B�7Q^�"@��h&�'��{OeY(�*��!��@/IRff�C<�V�v}�=��s�����G�^������ɓ��f���G:W��s�s�F��Ȳ30Z�9綈����.z����k��@�b��HN"���&�1������2���N��C���T�:tx���W׈}\+�t8�`"�s�9�e-.X[�;cHi�+�b�����;� >8�(xq"�A�V!��"B�YvΒ��O�S
���>h@3k��QJi���r�:�U4~xk�׽D���y>��%���eΜ�A�g�u�&�b�Clll�V��t�;w� �{���]�L�iVLo�?�?�ү�گ�����Y�)}�lr�f��mKfa�%�HH@�P���k���Z�[A��o]"���P/2z`�(m���Q�yo?f^R�����q�w���=���e�b D��B U��Xc�R��*Q"bD�/>HHB� A�D%�+k��W� +"�	�FR313)�t��e]�˺���b���K�}f/�Om����~���-dY���0�L����Z��
E�������o~3�~���Ʃ�-�������U���c]ҮÓ����Z��A�RXA'�����f���6�� "D�s�p|�:��p����C��6ډ��$ċ��z�ZnȐH�'B���\� 9 �&�q�ИN���i��b0��H O�!fM�}`kmduPꕣ-/ū
ߊbȂe�W�o��hI�ॗ����3��bVL���I�N��:�1
��֖ ��Q�=E�� p����_�tx���>}�;���Z� �L��D���L"� @���]T�����^Glj���*�{����ѣ�� �(����v���x����:Q��*}ǭۼ�>��<*�)��ޤM��"���dfx?.�:�13����i�I��:Q�;����V�ݼq�{�(�,� C�9sÍ>f��s��eQ!� �ij��A$yֻ�on������S������H�]f�ƀ��BbK ����zi���0F�V�4�6s,G_�:���Щ}:,���I�����!e-���z�!���2�h]Oo��kq.j�I[J�<�\�&� �M�D������S��E�/�p���}!,����^�G?�Q�>s����-����j_��V�$�h�&߶3��s�_��_�8^0<�;U���p`�@���wU�6D+�*Q��(Fb�# �߹���Б��G7�u�P����Y�t���f�ZYRט�ԫӴ�a����ץ4Rjq����Mۦe"��UU+h�s��]�~8�{0�ϑ�9^{�5|򓟄��,K�z=dY�;��6��eY �4y���*���a���W���~�N��/�������rG@v3���l2�['N�����c�q�rVS=�L�&AE��)�$���CQ�0f���:���YO���,���]m���y���GᨴG��[���A���<i�`y]*�G���qT��z><H�����쿣�J"�8�����p���W�պH�"V��8LZ�|�^�m>h�i�u��u�~�w��yy)�М|�Fa���������.�3`{{���'�$��[��N�:�O�=�d��O�������+ ��#|/��F��W_��ߟwtFw��ǟ��'gI����I�M�1���ꢬ��@�A���P�S�^�`�F��u�p0����A[�jGyv}�p� m�|9���"ǘ��1�ͺ1�<I�4�x<FQx問೟�,^}�"���
�~����p��M|���&�n���pk�Iʋ��w���_}�T��S�zU��׿n�^��Q��J���Y�5��ΖU1T�9I�*ɒ���&676�@��$�,�+��l���Y���?�>��C�Ԣ�9�A��p(��~{��6-��kCD�A��Df I4�"xo��p��ŋ���ckk!�z�y�<�#�{`����0�_*Q����n}�W�W���_������Lっw`���K(|;�^e�NΊY��e���I��Ι�8��^�\�qeY@)�T^p�r ]����z=��t<�ѣG�i��������|���w��1��qǿ�$�q�A���D��t�T��/MS�Ԧ����㻿����k���ad�<yŬBUY��E�߇��wG�����ɫ�;= �_����#�P�g�;5���'/��3+���~K��D�S���p!����>qr���Š߳��P��$�;�M'��"(X��=�*=ݓ�QX���t��}ʎ����3�(p�>k�O���,���I��У/�1�����>}�}������_��!��41M.�9�#��R��z��{8{�,>�����q���:����O�<	[9��3L�%��iT��wn��	�N��?���<Ҋtx���J� �dU��
W��/�$����_*f��^B�C�~n@Ӽ׳y��T�M^���B��#�S��v���Ӎ���G{�����yW��t�5�>(b�~���j���+}O����s�~��7/��(�,K�$	N�>�4Mq��&Ο?��/�ĉ �z=�GwB����: @�|�]��Z�����v��V��3�V� ���a*
C��>#���~os��^���Ui�W�$K|pN)�$���{���F��,ଅ��������ĕ��Mz�U��;��xԤ�Q�q��G���Z�8��o>z��1���?�wl?��w����~�m�z�u��A<Z366�8u�Μ9����x饳x饗����(ב��Z��ޞ�����1�ͤ��{U1����tK�u�궹z����f�u���KL��`�����])ڝ3"٪`�[;'w_��˷.����ڀQ�0����1��?�N���#��;��?G��q�5MSlnn⥗^��/�������`���[����{�5��)��@��ۓ$�RUe��J��i�X+����
� ��}�k��o���1�L&��A~{�u�����~p���������);33܉���IY$voJi�(�f���z!�JA��^����&��8�E&�A��񷸬�q�\wIBz�N���#\!����*���8��0��m�0_zx���܌"���:y�Į����L��`�.b2.���9ݻ��r���Ǆ�1--}��k�5eZ�?� (Z^��}|��,�g��Z���o;��#/�9�bu�����f[X^�`������i�X�+����o�w��ς����P�˺O�:�q��n���s����X)8���[*C<G\ybu\4�,�=��j~�����b�7k˥v_���a9G\���2O���i�a���v���	/ƈѦ3Dc�=�b�Z/�)��$3�97Oc�X2��p9��u�=�ݞ�_�� $	��:�X���`���^�Ͷ�9L�S����g�;}����!@��߁swo����;w��w���K�� r�����ކ���wn!�����7��ڿ����� }s�G>r#��>&����'v:�}��Ib�щ�TU���$Ku���ΓىS'�k�����[��;{�����H�(�.ԄB��-� GY�c�+ R$�x�ѫ�iy��ݣH�Q�����p��I;~_L��'�-�b����v��U�О��ui�#N8���`��UR����#��d0֩MW��&KXS����H-ױٳ��X�4����q�:Z�i�����'B�4�,��]�vߵ��>^麜���O�6��y������m]>��A$pRH͵��PUJ��9"Yr��2���r�:�T"�l6��I�W�r P���>\��Ƙf��v����kκ����H��X�Д�Y7c6���hD���oږ��c������6Z��<�Q�2'ζ�^݆59�~1fBX?�e�܂<���ً�ؼ|����곤��]��n�Y1��.q �e	�666���1�q��-h�������&v�<��    IDATv^�Ω���
�{cTU��~�����>�*XW"MS���e	�1�2���&|��݅s3����W�^�z�õ����a���i��+Z�[Je}R��U�4K�,K1&U�1��z`����o��y��M�g�z.���u�>�Y�b ���y �����	��t{�<G�"<���(�������Ԋr�S�:��������-�����:�����_|�o?�Wϵ��V")\/�	��}���M�"'���'����j�����
q�5�)�q���o�]�u���uM�޳�j�����:�6n+AD�(2qR�u���*Xk�$YCļ�ͲWq�6���eu�c��Q-�uH��9o[-��QJ�Z�(j�,�:���&6u,��F!���4M�k�[%=�ǵ���^��4MQ�%��+�r�R����W�U%�M���^%�]���.�s���?��mߧ�~���ƶ�Jg��C�����F���}�6nܸ�,�p��Yl�z�?^����Ac6��UƧ>�=x���B��_�1��0Q]g��G�L�(�+���c_�/_�r��O��>�?�]G�{��o��ܻ~H�4���$�����_����Y�J�P�4�3d���i�ʻ���$�~�����y�����G`�B A 0Dh!'��Ȃ�3/���C+u��v�x$ȡv��S�����C�C��=����X�.�0����ww�q�W a��|��U�\:��~���)_�:��z��X:_�	#�����C�˽�������^���������th��D��G�������3N��2ah����{�Z��������2��%"`�8vՌ�&>��B�{����@UUK�_]�UHD��)�2��<�6̲���&�J)h��Hk�L�~Q��n�+n/�r-Q��&�^:.֯m���5�Z����`�d
o�z�s���kױ����n�����S헠uc���^�V�G�g��g,@�[��v�m���R��~s�i�$�%�~��e���1�
a6��Zcju��*��H����}{��)�Α�H��Z����PFa4�C�ll `m���eU�t~oT��N�������]�rep�ʕ������w#�c��YQ|S��|Wk��^oP�keU��ͼcDBe+�����i��=,��2��
��1X1���� ��C�jӮ GġESp�[�:v��y|8�'���k>��$�i�A�r�vB��a�')�`���^<H����O�,�@,@ K@@ I�]���(���� �

Pj�vi�������b�W2(���Z,߽���O��������ʣ����Y#MR6p������= ͏����ܨ�/J���6ɉ ���.�H� W�Wz�\��=��:�*m���*��H��9vU��][�i��/~��#�J^Y��$�L��,��i���ܼ-V3/O�(��h�����KkmC�$iHO���~�~��,K8�`�bY�$I�r��G��LTۤ�.B�e�<�ֺ���~�'��J� Sm�����jz���{��������n�����)m�3�IDP�e���y�<�e��Z�5i�ĭ�OJ)�8qb��3^#�����%��_$���J)8琦9�,C0��*��N���� h4 �n�� ;;;�o��B��{{�U��V(K����7�����?�?_��?��3W~�J��u8K� \�tI�<��Zo���`#1C����D��%ȧ��,K%5�1������&�u{�w�ڻ��n��hei�� ��H�A��U�C˳������ e=6i��P���ں}�(���G�i��ïϭ��dd�\m��uXU����u��u��:����Y�t�գ���quP9��V��^�7��J�	��*Eј�V���sr��t��a�'�֪p��N	)��2�V���:ڪu��M��HE��d��H�VդU��n�6I0Ơ,KE��O,�lV�إi�,��~o��\�d��Z'�WPS{�KhaN���sB �f�z�}h��,g(�
֖71� B�N��sq~=�*$I�$� �9�RcR������) !Ծ�����'���5��ޣ,K��(����Hh�ב������8����'c�y���m����j�|-�tF"I�Rf���9�b&�K�d�'ܐ�<���a��Y[5��K�m�m���	���}3�"�t�5�3�e��aC򫪪I>���y���w���7Bo���g���y�&n߽��(`�T�w����A�o�������_)�\��[W��ӻ�@:��PIP���3��l03'M��։V��}�W���<K��r.��i/�43 e��8�v�;��w����=�2�I� F�F3/���Q�*�Q��ㄠ��2�}|������"�>�?�|G��z�<h.7�N�h>�������7��'���Ѫ?�:��J�ڦ��b�6�����b����?P����0����^����>�ܹ��h��H�&4͹ԲIk����fR^%�"�4S�
���U��6�j�'N��l����T��6o�rEu�MҢ�U�H6"��L&�m������ �nUU�iq0`8΃K����F4�NU�V�r(60�Bb2$��V��BeKx`]	g������E9�b�43�����3i8W�*\�`t
m����MK�`a�<u+�I�Um�$�_
˪� ��su ��<�/<�C��G�1޳Z�#P% ��h9� ��i���~T(��h������Z�,� |�͘Q+A@��*��j�Z���.�����X��A�1��<�c�Q?�����ss�n嶙����gM����m3'�u��֪��c��������t�ɴ�d2���&�Ҽ���mܹ�k+y�����`��~�O�/~��~nt�C�C���I_<�������O���W�~f�+x��!ȧ}e_~��A9����:�]A������}�=��aooB\��5~}��F���aJ�B��Z��P��}�v�O\�T�'O'=G�(��0�t?8�x}��YM����S�$�e��k�LŴ��iژ�bPF|��f���Gr����|I9l�mSO�H�	b��_"k��ŋ"��<jD����qRUJ��YS�U2֮�AJ�`�[�O������گM�������?˲l�Ik<gUU͟���`���~��O�UUa:�b:�6�9�&)'N�X2oF�e5�&��H6b����`{L���n�]����Idiִ�BiT�/>��Q��D��c6�-)�JŔ/u4�IL��&��s�9�9)��Y)ds����x	2'm����$s���n�f������Q�Fǀ�,��=�R & ���ʞֵK���KY���sEQ��k�8c@2�Q��8�G�@X(�޻:�̼O���b�<��4m^ʪ�p0��j��E��e�,�1>/b�͊1��:TU�J+mS���צ^ ��_Y���Y�������Y����ǰ��N�;ބ�B�����2��5��+��g����>D;tX��"} �˗/��D��>m�R�n��}��R�7�?jg�~���y���i��F�Ėnp����ƍ박ŭ�w0�`t
cR� �a��h�m��ќQ��'0F`��U��c<n�S)��1�ALC�����SќI�RY��H�=�B���n5o��r����f�iO�q"��/�!��=�k��o|�����b�g�T4�O��`6�5���(�E$8q�h�h�����v�^u$oO���%B�$	��>Ҵ�o�6FD�B���&�<�s�Q�vvv@D�lM,�/Sl��O$h��i�6�p8���.��h&���Փ4M�RUU=���7f��p�`L=���]���X�����4M�mj���� x���`&��cL������ʲ|~�rZ�����B��&�跴��ь���Y��r�ǣ���|E����Z~\2W^� �^��c���e�2�n�:[�c�/����{Hu=>!��=�E�F�Ў�m�x�R�y��o1��DP���CL�R���ǘH�3�&��eH�UY�:���<R�ZL�$&i귪�:��$�ι)�&����xi���\��u�������9�<���	��s�u>�P�~�ߐ0V�o���
A��?h},"��A "�����O�⠈-)� �>Q�E�v�(TUiʪ�B���AC�� @���QPJ��B�i�".�(��t[�V� ��%`�"h4�U &��V�����?��~.�O�. ���Ν�鷾�.��r��+��x:�_ �M<��}g����/�ߡ�x��/^��_�rz��;����`��OhCQn�E":����r���Z��t�1͒�x�U�0OQ��Y��x��N0�0)h�@`�5�Q���	 +��	L�!XW�*-�^V+���<$� ��P���i�7�j�@[-h+�A���1�����;$f��,�1?�z�F��>Ey�7�0^?��C�e9Z5q�	fkk�1_E�,��#�&����s��lS�?����S$s1:��NTVΕ�5�iH�s��%I�y^����	3*M1��s��h������M��bT��|T��m'�8�Gu=/�}!���X��9�D��M-�M������*g����TB���OE��&+����T�t�U4�IӶ렍��,ʲ�u��'��/�[�H{ۗ/��2˶�p��+�;�2�Ib�D�67�y�a�J^$V����aE��"��W.��]z���lU�HA)��F����0�`���#��|=�����C�j�"�B�9�����_<��������ypZ��jk����ֆAP�}]��Kkh�ʲ�1	B��y"q�	�X�֋��Ԗ'�� !	B�P���&ˊ"DD���@$�a9�IZ�Ê�3��z@>t�\����xϹ��x 4��$}+R�BX�E�,�$RJQ����2O K �CL��9��'�@`""�P�EH <�aR ���zAsP�,+vD��k�l! $̐���$��I��;@"A��B">!b�U�+b��Y��_��	#d��UT��t����ݟ��y>���?�L����A�  �/_N�a��]�PN��O���*����dF��aY���a�;߳�K�,�$�Nz�0��BH����N�X�QUD�(�i�<O6cR� B����ij�ۊ^�,��A�h�icTs�Z1\�����تI�p8�p8D�e9��"����⧔�x<�p8D����d2i�^���<:����l6����� ��d>��n^��R��ͣ����s��\�:|��R����a�##�"M3��1�ჯ#���H �4C�&K�l0)H��6�B�#&dUK�.��AԘ�j�!����è�(�k3�yZ�������o㱝#��j[��8��<k �s��E�uDg�Ӹ � ��R�pE�)��lND#q��D9��s�U��¼��m�w�?S��ڼ��^ӿ�����IUU��!oT�73; ,�T)^'�+�l�JIT�j�#�I���/�H2�@��+"��M~��פO� "�+�zH�E��9�HC)��0����yP�dA�h�l]pD��5�@��H�/����L�&B^���y�l!^+dV����}W@,
�"u�w�y�uU��^o���nN�4���LJD�H@�S� �'"$@��Je-��*[��2-�����	@��J��r�tU@��HB�E�D��G�1���H $�A�AAI @������2 ���sW,AẀx�V|W@=fQB<��D��$x�����)	 1	D��f"�~�pD` 3�ibė�kbH^)eCDLM�������(2b�)E�$�'&H1Dd"H�2�� U�{K�f���Ay	��#;�wn��N7�����L���G60��ߴ �ʕ+-/�>��7��{��{�0εҼٓ�U����T��,M�D�t��̺��?���;�ub��^� M�4�$�xv�Bو�H��677[*��RSTc�!�m,"jT�����Of�[2��sE�0�����H��&f����*���P�A��2J��%�|���H���KD�Ρ�*�������D�Jկ�<w쟓�:��CzC�S:4�~B��O$ޕH��A��{("�୅���5Rc�ZCs��! I3���ے$�u����{ddfݺ�MQFR�L����ؼ���K��z�٘���Jf$!U7Ш��k�����<����F�6���~9~��s����:�k,�U��)i	��{kG�UCeA0���9X� T�bɵ��&$3�8>�Ja%�2b�,_��^ � n�w�5в���-^�V�(�c�r �����Xs��3� ���{@+e:^gS��cV	���%�@�(ux�Zz���������ܘ���P[�}fh$����C��df$�0zD$]\\�܋��{I� `�,�ٶȔ��ڳz��<"Aw7���� ia�7my`�̨��XI���ԡ��Q3��Zދp�ʵ�#	�^m�������$ #@3/f�$�H��+uiXҸJb*I���c����X� 
@���5��v���2�e$�$4��w ʁ]2�sl�"C�Z)H������&�d$W	��=�Rmm	�F�E���g��$�@l�F	� pA}>��/ R�(���W�JZ�4��\�'$I�z-�nM�[�f)K'�p'�F2�S* D1 ����ک�m%xEr���&��##/(�'��mD��v&܂hi6��2q��%6 ��-�-V��kt2E��EDTAFh��b�w�j����=i+i"�vfv'��H�+�Y�h�����>��s���m������=�����������������O����T�e�9x�ʟn�G�/ß�c�'�0���l{r���N��R�����0_G}�a���uj鬐����k$2���� ��������G'���������]��a��~z��&6<H����<ߧ�: 뚫u] �#=߽��>������S�=J�?�ൃ�^ŷ�4Tv���NN6�˕�7N2�`�۲f�^(�nΖ�S	'n��ܐh	��B
�XriZ�h�i�D�� ��2-
����ѐD�	�U)�Ī�(Kw�4YA��&W��2B-!+0�2E��.3�����s F�$��2	�18��~��Ps:�fT�L��*�#�be)d��0���`BA�a����v���PI�̤����T�

4)�L��f㍹M]H�$P�)d��L/t/���%Pf�D���%�$#��,�~��\�2QA�R�^��(QS�H+���֖u2c�֧��@�P���}D��RH �G�	�_� 
JI��!#���:=Y n���}�v���Ğ�
��d鳼1"rE`�TI�)�h-/I��l�@b�
Ҁ0�М3cf���A ��2@ �4���3��h��o3�k*�F�SP����#���f��I�+tC/���u����+�@fJ���L)�H���QIb�q$A;%WAň!%8�;A'�m��  ��J��_)�KȾU�^���NED�7	�X�k +�'�8�l����=I'���6�k
��4'�Hy �m"�A��ɜ� ��p-��M�yVk��T#���nU �������ni �B��|&F�% M�`Or��IR��%��?북_��~�ܜ��'O������8��c�>���իW�����G���N�yi�+���"�|���T��t7e�Z�l�O`�֩�@�2ġ����x9�O���qdɎ�s>AB�p�Bz�f"p�jzT��ʠݛ�>�a���M��B�h�;�6��8s�������t�?4�P�5��.�D���H+�Yk)���$��Q��3�\���H){>O�{�ہ�."=�v �Q��)$�v�9�6�	 ��F�aZ铨g��Y�3����0M�v�XB2t�8����L;��׵���Ief�gt�X)����������}vP3�sg�jdP�Q�%47[����1�B]�Y{>-S�'�  �IDATϻ� �2R�y��Պ���80:<|�gEĆ]`�#���fB�}R �IY�$.��P ��́��X[�� 2W�Q	,��8Q$Ԛ��_�֚�e���fՌ�nT��[�sR�ݥԤ8egD 1��"A�1��,)A������3,(JU�$o�>$��=2�Hj{�5�M����Ho� �a��!�*�$�9�	��-�;�/��OI�SZ	��䒉;%�ILNlEn��H�S3���]n3󝄕�		�TK�#һ)H6�n���Dx���^]j��!͈�Ɔ�J�(ak�H����"?��-3�B�h Q%��ߴ��ɖ�7� �L���r�\�]�E�B�Uٞtɥ"3P%x,�=��@��V⍓�('U��q�d�RH����+��{����Lc"E��\͆�\���U�G08����6Rq5�F�3$�L�-�&���*�+w4)���IM��t�w�ߺ#����$2�-���5�朴pG��(�� k-�k�gt�TgH3����Ӭq���f���&NOO�f�������_��o��W�^�v;��x���g}@�Ꝧi�L_���6?����/�C/+��n����M@������8��$Ǻ)uܞ�T��m;h,�����=�8�����ﰎ���x��#�Ɍ#���*/�;�΁G �R��(�`5ph;#C���PD�A-"��A�:�$W7��-��Ks�=���*)�fls�w��T�c囓M`-^n���m$�������m�k��[@��F"�|]��B2(�P�d��3�b�������ڕEY�|�wo�͙���s��O?W�g@:�4Zs�5�W������L܁E�H- �N��WI)E�Ҋ�eY���.J�p۠���!` 8+u����	��n [6�͔�kk�����( ���x5)��x#q6b�Y"e,�˺�wo���,<!yzD����~�����ȑ�9����ImP�+	; ��!'�čB3L����aߦ�Nfb/a!1H�i�:�`�"�k�)�f0/��~��Z���'f��r�S�l0�Q��s O��g����T~f�gF�0�.�k�R�\��݀�!ٔZ�^Hy��i����e���� .����f5	�������ߍ�˔�ؙ1$EH�D
L-���vR����H��B�!�s	{$/�!I5�A�.�?P h�0K��( '$nIJ�(J$�0H��n�_"4���쓐S�D�<S�U�Ud �A@��um��+���\H*"7f~����R*;;�R�LH�6������d�_|�/hȬh�$Z��R0�h ,��KDld\���v�kF��b�j�Q�eb|)Е���
V4d{Lyr�zY���� r���8��` �%w�1ǛKRb���ZaZ��5
IX+���4�P_Yï2��L{W+�Rָ����zJ��lssz���;ȯ��*�����=�w�ޭ_}����k�믾�˯��C_8]�����_���o�����������_�ի�����-��|����EU��,��Z��0�i�4����8�G�mj����A�r"Pͬ���D�ѕ �g���, ~H�t	��;i($�~�F��9�\�eCGx7� �M�i.���  G%52Iq��ݲ\oo�-3��:b�1��p�S�F#�&��*����\�y/7F�N����IO133it4�\D���)!�{�M 2%3���fZ�"��г��֊�p�EȚ絖��g���\� ;�� ��s#��0���?���[Y��; 3L���\��d��-:��.h�0)���7����D~"� `�]�R#�~a��M�|
�3 ��ncm����	����w�~���1��k�3|������ߓ� ��ไ3
��wmk��.)�q߱%�g����i��c^�<!��]&tA����[C���F��F�fƧ��<Д���_�"��(��� |�@�X  �[%6N�*�6�.�$h� �=]��,�3 �J���[#/	m�)��4�)��ĵ�Sx�^{P%�;�{�F	���m�.�ې(i�-0p� �� }���L��4dg^nL����܆�"�&����r͑կ�r�(&��y��%�;I7�o�	if����\R��D3�-+�%z� '@[4��#y��}E�ȬP���wsY��G�Ӣz��f.w�����Z Jq钭A`�{� @�=؈@9� 9e� d:k�{[@k!��� �sRՒ3
��C��Y���-�e:��<���V�/(xZ��F,c�=��Xչ�7f*)T�eڍ��L|6���ʥ*��lD�(k��������>�Э����͛�>xSk\����Zk��� �Ln�Z��,w���`!� �Oc�ئi����NNv����z��J��>׻��ś/�͗��իW�c�������} �ӟ�����nj�'������l*�_M�|�����?+�gn^H�����͆�1���Jq7�.����5���I��3�� ��@�vR��� *�VX%5��A��4)�̱��W;�+׌Ʉz֘G/+	2�F�5���ܴ�g��ˌ8����R:3c�|ۢ���)�Y�&h t�n�ì������V�$9�B��.�fU�W7��Z��P�@��:��eYwkks��9i3�k���^~'e4(�	��כ�Dg$�م�B�R�m��	If�
�Kwvyf�8%���N`lۥtr�� �EK�]223�Pb��zrL2���R˥�C�ŀ�T.���v��D~"�ԀJC�~)7�)u�J��h��%]��IFP��Ab�sr�����$]>��� 3䚀���� ��Ժ��^�|U�%8#1��B��̼7)�N���a�zuHK�c�dy�	��.�*��	W����Z �t�@k0yxfJit }�?�?l��g 0v�%ݍRKX~fBK��akB�H	)�M��Q�Z��_����B܃��F�P&ҽ�݅�ѫ�#Jos���M��R6���um�R�ko+9M�L�<��@����k}��w�����e�p��_ʬRF��MS���� ��d���q�I�vw�ֺnطO��|�u��~��N����z2 �ݨ�:�o?��D%BelH�-����C������,�M �>��0WL��^�]U���YK���sؕ��~�eZƉ�ɾ�����%�' �a��4ޞ�v����[�8��
 �6��n�?�=����˟<�����ܞ�ɓg�!߼�B_~��^��J/_~�������c<�s�AAЭ\���FI�M��fu�/	~2��8����?+4V>#����W��҉f�&���TƗƣP;$n(�ӱ5b��LI����7�HQ`V/�(R *�eu��g����dH�h&5>K��id��t�����
3��NK	��B�����
p��0W�S�߈�4�M�U H����m�� \�-�u���J����q;όZ��kD\R�IF�>y��-���Z!5��D*$:��)0� @E�3�mf�+RA���$M�}s[{i%uH�5E&��x� 3����DO�Q�" `�`�,�0�JQf�J���
q%R;�H{ �������$��0��0i&	���̔��y�����L�d�(�/#��.����.-���(�@���i��?����Z���³�x�̜N׃֨�r`g#��l�ZoKQ!}<XY`YZ��eo-�����E���a ��{���,�e9M0��Y}y�o;��'����uX+[��� \�8p]g�:>Lo0σ��;��p]��6��eYUʠy^u�G뺰��q\8ϫ��է�O�5 ,֥!.�fX�}[�ۍ?8��k?����у��:}��|�߾̇��>^qh��ǫu�a�t{ sð�_�,���3w�u/,}�����q\�����_���z��<m�������.���۫~-oa�ߟf٬3�s��f�A�����(Ĳm������ v��w��x��W?xN/_~}��ի���6� �1��?8��W�����o���nv�� `:�k��,���3񒴉�k�Of�A�_�`@R֋1��=L/�Lu��ƍQ/H���{�P�&�)�\�͸d�dC��� �������U�p?�Y$VB�LUR��AO?1�i�ש|����h��{ !r0 �v�c���4ebDv�����(����1���=]�v��,LLh�AQ$Y�7�|XVZ63Xʰ����_m�h����|5++�A�d>e�T�<3��ߊ+���d+��%�V@rgƝ�-i��ꆖ�Fz�֙(��,ꂺ"�6�`fm�0��j�)V_�դ��=f#
V���'w�hfvkV@������fV#su	�Ze�ȭ�uW�����꺟5�Z�=�N#����6�~Ts�Ojp�c2�NO�ED��:�v�SEo�>׋����o���>\w\���;}��x��+�˗_�͛/���� 8nw\����a�����_����V p~��wi���i����xr�A�<�	<�8���7�{NS_/1�a���S��ސ��Jv��ZƱ��c�����wG 8Y>�P�f�q7�=:�o�z`7��$�ۉ�2r��sYfN��;��$���fk��i��z���V纹)yz����������|�m?γgo���}�;��O?}��	h~�K���ׁ��?�^�ze���ן�>��9�����5��_�����_���Y���>���1�)����c��V��4�7c7>}��_��!�3酴�3.���XO�� %�ޘC0 TB'�vNh��7���[*�tG�^����L��>�N�>�&F��pD&�P���mY��g���,׶<s��B�+ɯK��� ��xY����\�J#'4ݑXH�\[�@�j�[3�0r=T�Z�Յ�ȴ-����P�����9�8	��3|=d��^�e���ζ�"���
��b��a��E���R�KQ)m�`�9Pb]�܋�|�2oUc�[����<�P�ڙ��� �8�pW
��K,�iXі�2�h��ke����9�$����\d5n�Ǫ�o�Lӓ��g�a��cĊ���E;?ǰߣ��5����\Ob�R�6Sm�5y9_\<���Rʙٮ����N?\��!�t O_�9�ޯ?=,��^
���k�3#o�>���#�:h�7o�����_~������a[�3'�u��x/_~͇�>\��s=�{m��7��9�`��/�!^~�/.��˗_��GV���ա/� �1��4����O^ճ�����~:n��$_��!����2]��O;��Mf�@�!qE`1+����^�]| �J����N�v�׊�V�j�½�k�rH��)��c.<JA�>V3���<�}�2r&=��x+"[]��W��*��e.�e�(�ԝ�<_m�mm�4�-��,eЪv>Ȃ6S��tW�ڗEcC)�J'�9xk�9֕��4u��a�0�˲�f�����Z���C��I�]����q�����,�L;%�%�\{?����9PV2^�Xݹ������n��2&�I �d���6��%6��X�^e�s4�~�+e_���f����,���F������v�Dggo��_�;�����<����}��>\��I���#�x��x��x��o���> ҽ[��ۡ0W/n���h+[8�+q��iC��Zc�CT.�ʗ���G�0���B����S>%=2s��P�P<5(s�b��t�iLN�g��+�Ĝ�����Z�s[�7m��c�
 eַ1�S�=���|�7�� ���0����nW[[��C�J���t_jD��Ϙ�%:��o ���M��#�u7jwW�r��"�g�%�m��ۃ��+Ǯ!��>��`��lnm���!��A� gg�����_�`��__�_�I����<���x��x����s�Q��C�?�i��ؖir��l��"���Ɓe�lM��>�q��u�6 �����ף 9[���ib���RV�y��\� ��]�W��Y�Png-ۑ�Ǝ1�4H��q�C��~ G��t���@tqq����_<�A�c ��{�ꌞ=����~��y�+ �?}���<Ԁ�P|���ݴ>���1�1�1�̠�a�'?��}��%?}�������/~L|~�����ы.>{�#ktd��/���x�� �~&����~3XzD�����������B��K��    IEND�B`�PK   }Q�T��!�D�  Ԟ  /   images/cf2dd1a8-295d-437f-92b8-7fcc138ae9be.png4�uTT]Ň��z�iF���n���n���)���fH���|k�e��̜{������މRQ��zM�a��J�?c��4�<u��Ar�b^�+]޹��<�B{�������\�K�B�EБZQq��SH�y����87�����o����b_�,��9X]�'�O!_�YM�cMO�S�ր���nS�[#~'���SB{��7���	"ݚ�g��)L ŪU4y�����[h! d޽�v�YHl��T|�S�F�>,��	�Qr�4Y�@>�T`Kc򆓓3�����=<�$$$�?�dff�°Ȧm�A�\W4�^l��r��!S%u��m�=�-Uv�q���)$%�_k8���恢�u�����G�j!��A�(g��r/���n���OOO��\�H�ژW��}���!�A���b�ԟ�! �0�,~*<V�i$o���=_���YD!�rL�ӶyV6�y�Q��>�K;�MV�+v�3�0-���c'1�] %x��8��������.F�6N�6�j����N����L��z���D�u�����ဂ�Kh�#�R������۴Ϝ����Q�J�w5�'�TB�G�琄����q��|����ٞ\9�s�\Ԟ���A�AEA��s ��Z5���͟���<s�P��I�̋�ƥT3�Xq���fFZ��d�F�h錓��Y]����A��ur�bR�n�쐝(�0X<(a#���Ό��Zg30�2dq���ai֭��N�\B�p��n���M�ɴj��$"Tޥs@�a}���(�B�3�����@T䘘����gs�@?J+�&�4��@~a.��au��E6���"�s���s���-���u�n���b�g3d����L@z���L�͑�숀r�{��͇5ua��p�����52�)���~I�ό��N�x~,����TI$qɁm���>��,�4��_:��8Ej,�nT,�"�dr�3���zmj��(>�>5Z�7�}KK��,��y��U}�8�d�ݝC	?�3U�9�O��}&��̬,1�n4J�Ŧ 
`	uk���%��#Ȟg�� q3�(Q��> -q�:���Gq���9����A`��QG,.I&���Y��I@b�����]鶟W~^
��a�����O�	�镏�~��2Ţ��;��������/}���;\���-8f��v���0���������U�4�;d�U���h�OK����L�/݈_��)N�"�'��!N��sFr���i)�i9���I@�@���5�8�ۈ�|*;	ѝ`0M*hڂ�PNX������M�Is���N�����a}�������ڞ�(�����`�5���X��هl|��2v���N�feC
R靾,�X�d���b�J�>A``�����Q�F��=)f5�������kd�3?*|c�3��!��(d�(d���Y�"c��2�����W3N�+�Ӻ��􆇯�)WZ2��حwSt�n�`��
��u�&)W�a5/�#�� �xз���۴ח�_!��y�g)�n�������GC�I��qԨy?�ZS�WB�R�ꝓ$�{!X�.��:F�!nn��Pξ�Gbl$V��+����N}��N}_�P_��Ȩ66{�ZO6�W���J�GMmm_�I#��ˤ,UJ�W/b�I�YRx��~UG�u_�6���,�wan�ɔ�2jŢC��D(O���;]$!���Or3��.u9�./���=�[��u�^'-�6T��D�?�x~��H�/;;j���5�R,M��ݵ/�	2����"7�掆�G�M��}gI�j���1m�l������m�#����|��K S��JJ����tV�fqZ��f��<{�x�{�o�D.%k��76�Ag�LD1_Y0�ˋ�j�eP�8GCVqY�0�!�o��o��9��d(����YU�s]�tY�~üxB+o��U'~(<}8��zN�\�a���1
�ơ\l�_���4��N0�Z��p_-Y��Oe�m�/}��2L��6e�N������}7�|�v1�m&խC��|0��EI>�"�j�6u3�B�[��p��� ��F�G��AB��w80@�^K��;�Z�g�K��_n�$ɾ�qӭ��1i���������$HL։�� �#�,2F�F�	$�8CB@���ʧ*�q���G{j2L�UZ'A�����ۏ��=��m���Ï
�o�>�XB�����q��k��K�h��e�`�aэ�ܲ�3�` =�� �"��օ��������T�lwq��T�l�,.��h��樻,�?>�?Q1���Ԙ J�bvjD���i	�$�������Ӓy[�4y9��Ye�����
����nad���;o�(80qF��� :�c�ǁ�YN"7�ƣ���o*�ߚ��"EyQ07�=�Gb͏�dc�g�3��gB'�LJ�K������W���͚�46
&��H�Dwp�}���R��{+<����,9������݆W?>��p	�š\4BH�C�83�#�\�a(fP�8t')O�3Fn�t�����n�H;.|�uE�P*ư�v�Wn#CV}�PoΩ�	Ҫ7dm ?��"��4����yV��ʊ�$UH��S*j�lWM?Դ�l�V.���]]]�yyR�I�%3@T��<�P3��c2z�BN>8:*{%�{��8������YU���N�twƞ�u��9j�c�{�t��B�ȑ-\J�1�60��7Ev�O�rgreS�$ޤ�I�"�����SZI���B�U-�ۚW?�ʱk��l��lD_po�� ʹ�q�ܔ�~�J�NCo��8��!x�Z�,Ftϧ��̜��h�w`M�������"�uT��ONmB�����gm�Qx���L�c'�\>����Qt�7�[�\�MH6V^��Y0Cq
���a�/���F�4a���B��6�jX�پWTV��\��4Z/\���p�*�r���sѬ�$�u2>��9_D�mp�M	��P���hgc��QS�u�kӍU�;�
ի)Ra�d��ۮ^8�n����7�b�L
�jL�N��x�Q��{����5��*�>��M�����oEҠ�i�T�%#&V~�T�ږ$O�m��H,��`�z��;ޙ$=�~x��g+���ill4�-2�Wx+���ǲE��~�#m��co�E,���T�jo�v�xa�#WWW�E��;��yX���ԝD��Xo�Ir[w�ղy�g�V-Kjڶ�:�܂�Yy*c�9�T���	G�����gFI��B��+";�I���ݳ����u�I���������|Y����(�ꆎ�Xl��c�gvU����v�90�~�V��5�X]��)f� ����l����pP����rwK�U�,x�J�}Tse)N\�2L�n��7�m�&�z5ZE@6 b �dc:�/d%u��C�,���f �$'s�<O��-x>??�Ƞz1J��"q�L�/
���r�Vl�X�E�zÐ�3����@�1��e�H׶C�
�R�G����]���z��$��rgٱ�n����I��^"���,B������~�R��x�rʲ�'����.���Ѝ�#+����՞,K�A����G
��pԪX�aE����4�mH�w�o�Wݴ"~x�s��Y�Խ3Q�[[�Ve��G2��-^L	��C�i��Th��<ʜ�zl�_��B�[�+�A�������}�i�$���
d�� ���>l>���$��)muj0�lG�������i\
�������%��.�]N�c0��	��S�-(���"������hHj�i�4s��8}Sb�<���R{I�%�&66m�8!Y��������MoJ��a��Y����X�覤�X��n�Cpmu���r�m�]B��=�}.�$�U��!502 a�Z5�R�uf@�L��0*�F�q�����[�$bmqm׬`���ǳlrّWTR�sb&u�,0߀�C�C
�q���}���(��y�G���[حu�X�{3P�qzS��8�O��&$ܰ�Rb��ȗ�p`r��Dȗ!��O�{�#�?[ф��l�ޣ0�s���z:#m����*e��pl�����)ӥ����'f�|BT>�e�7�a}��w�}������ԉ���*�;��N��R rOU7���X�Z�,-�6z����2ބ�-,���̫�jq���7�iR��֦7�����_�D���[3���6���!�73�P02�������|}�u
�!v��c�[1��E����?{2ϻ3S��w~�@�f�8g��*[p
~�?���	�:g�n=����)���xj��,�p� ;�ɳ�����_����MS � -Kq�=7��Ѩ�߫y��vk�
)bl��u��y�����Yh���WL�5]��%"Tp-��7�z���,�m��W��^^�_�	N�PS�*4���U��X��m�FG�95�Ь�̐2�	/
��.0�vZ`le�-�I���y��p\Qυ�2&��0tt�1#1��i�C�(�/��ю�W���J���F�>�"�4�_��L��T����i�f#w�&��ۨ�$[ɪe�;�W�(Skӗ{QP�2�S�?ł��X�]bz�Dn��;�,�L1�~0+��h0��F�/�k��qw�,摫�Jj������P��*���o]F�2�V7ց>3_Nௗ�N��"��g()�*\�>��J�SG0���H�v!I�Eg;�I>DQ�bn�Ji��!Ku���Y�d������j���D�s�@�̡��~Ϝ�/ԭ���B��>��~��U$|�r� f��G6��`����_Z�%9�ے��Z54o�Lc��,��8F����@�ov�kڍ���}�n�7bV�]ˈ��u�I�$�_V.��*�B����/�3��aL�,�c�g�y�[��^U�?��ـ���t����6b�C~Rb\L 2���
��`zc��~p�A>�V��C��W�}1:,M��V���y�=H���B',�Qm&�V�{qWCB9�T�Y3D0����ӈ��ٖ�,�:���S9�hW�J��`�P����;�T�}��6�3<��"���,�s��X����j�*Q$E���6�(�#m��3�f�.>ॅV�>x]�z��>UT�6�c�C��Q�錉"ެ�]�I�CCLVF��"������l|$���C�_W�?dj�.<��t-�:j�g��qde���;�
�ߑRŅ
�h�T 㸓C��ڸ��>�]N5l�S��d�����˲��D�٨[��?H�h�_>���V*H��h��u��p�u9��ˇ:��fT�E����Qh�^�/v���0�H��1��=R&��h̦¨�0���ƿ�0$�/�*�)QUj�}���ivZ$gި�	/��0G9{��3�Ӎ�@�T�Ҕ�������H�F�|g� \��-�kA=xl�kh�<�],�C��6\$O�n��j���!�U� :Z� Nx���ǜ~�Q��^�4GiAJ��h�<��`$����34d��-l@�6~U�+�|�b��Η�7��/s��3�,��;=e��\��@ 0��;���H�8dRh
.��ؚ5�6�Vr�D<�n&E�%OR0E|��o��y(�q�~��d���B�xm��[�,ܤ܎CB"Ȍ��==�����gDo
�"��q��]VqrX�֎y�����Fr�?ڒb�>�[�\��*���WK�~H�Ҙ������^�{�K��px�	��V�5�
�W	CN�YVb���t=S�Ϯ�i�1���F/>�[���	��f/Oh�r��ʈ�������i��oQ�;�x���yi���o��f���L�ypှ�ǊS���[��T���u8���fAp:�����I?vTj5�V���~�T0xM����{�I6TE�me���0v�z#g�I�ʟO�GȻ�R9�Ҭ��Q�Ar��Kť-wF[@��6Q �#CQ�s�"A�a園�ȅ63�z�(�S�u� ��h������7���x#����f�,� p�Ug���7�J+L��TGD7�b˟���N14� �����:�\BQ7���C2��C��c~�����ɯ�V�Z�>�g�X	��A��4J�Am۷����Q���/���A�gӶ �a�On>�A��8������ny�WhT��w8%����IC��D��0�	<��tt�`�<�.���/\WoF���|y̭��t�d��V��]���w!O#<�o�]
4�Iuί��oP&@��l��[|U�=�C�*�z^;�Kժ� �H"m[��l����5����M�o>݇����_��� ����P��c/������Gk�0re&�+?��4�` �զǮ�+��0�ơ������[�Pl�oR�b��i��Y�Z,����Zy��tqE�F2�tvâ ���R!3�@�5^{Vt�4D��^�̭̇s�����6����W�6�k����]c��A��q'F�>��-�K�ul�F��?��C���v�R�J�ίVE�U����Y�/��s�����$@,N����`�O����Ԩ��uG췖Q;�#�SңM
������&��fK��V�=��u���`&;����/��~zSV=%ʊ�=���'E~;���͚(�e��b��~���ћ<�<��Ej����йj�c۲��ݡ/;�g`�����6��ӧ�i�h
�<^pe���$!7�`�ē'��\[3�4����5ۦ�7������[�k]gIL���l��K�v͂O�C#���!^�BN��pAB��s.���ky��y�Jf��������.Eƍ�%'�m�$���7f�}7��^�w((>O>�-�!��Wa�L6"�(���f����%i�D�$W���K��Č�z��L礊�КW�Eˣz��x�P�\%���·}᭝�8%L����~L�6����u�{=�XE���NiႏJJJ; ���7��'�����-d��x�����?��۝K�����]{>TP=oܤ��Qx����q��a�<���|[��?�ӵ��?b93Zx��T�I]��b���뺊�oaL���#2�q�E�ޅP���Ý6-26o�bF
�}�:/&C��\}Uz��3n�P܄�7)�Zt�u�e���Ĩ��]Hw�P��r�����;N'm{�g�2�/�k�Z����L�(<O��(�8�׎�mOX˭���ej3j��]��:r�.������?82X0�^Q��د%���Q+����G���x����c������탊CכUO��Ӯ�gU _i��WV>�F��l��N#V��#�W#��3��X��y*�U�KWi�7�JX����V.��\�j�bj�I��ˑww�PR,���
 ��o�|�w���\�\�E���x#F��q����<g͕��;X�`uQ��^��T��������g�C���nTO3TO��-L7�K߆^q�u����k�����z�G�n???�Ӎ^u::��aн��g�	ɎN^t�>�k�a�҂���'���U����cS#%" ٥/��*�$x�/���2�T=�۪:҉�����L�����zv,؇��:�nV����_�c�����atA�YKF2�4^l���!xN����RK�� ��V��gHA���Z��)�9�^� w�1�\�ы��[;:b�8TTV6��!���*'��eu=��h��ei�?=�1�8�K�������s&���AY�҂���F�N�� �����k_�K�]���˭�{޲�L��c¡�=��	Dzy��b̖-#�RJ0�j��z�:L՚���]:�Z��>�8����0�~�ˍZAp���kIL��D��j4������9V~��/��NWEEE��t���ԩ)ڴ�h��Ԉt�+~�=9y�ofVV��/�a�$��pIf�)�	KNA�ؽ�@�֧��u�����#~�^obC�s����U~���2O:���f�����W����w������[�˭"S{;�'��z2K\�I�z�u�ф�p��I7Fmn�x���_�U��~(����ϕ��*��U;�*�B'��i�i�E�K˱5~�ZD ��(��?�U%W�T��_������d ��gj�P�!N�D0
��&���`!|Qͯ��a���
�k7��'�"�1��!H�2��殓c0��>Iv�]��+Č]Xk]*��ciɇ��h�  0�g~�� ����J���{E�lf@�4�"���� I��4Y��=�V�F}������>5�Р=F��k�P���	Qj�ZC����� u�m:�����4��������˔&�D�q�s����G�{];	,�q��:����Q��C�Z�s��狗�&����h����CF�+���xO�l'��;MN�l��jq��<�W�!��H�Kf��ݥZ&���0qpƧ���S����a�m�;?J :��n9�p!���dj���/K7.�**O�����"F^���%95%�>�ET�t�.|@��v0���F;\�w��P"��tn�v���"Ly���s���.��%���^r�伐D;���5j.~�9���Ͻ�~�j�Ȗ�e��J� ��J�e\D*&��Q�d��-�c�о��B�� ZQ�K�I���
�4�e)�466=����
���� �+��Eժ7�1m����8��j���Pt�= ��>�`�r��e�bgʵ�kO�9�|�_�T+��&D�͟��Ω�[p�W�E,�<�K�37W��8��)ˑ�L#���lK��7�-��h���_�~~��GIôU�L�e�:�>��b��E���6@��=^�dN{]�0��O)?��'��c?�Н ��Iy}��� Иf�D��ԉCDE�7����
%pv��P]�/�X�4=^���?���K���4,�����]2T������TH�y5~���F��B��Ae�O��w+åMX��/���"48�$�E���*V|�F�'#̮Z&z������i�Q�\o5��<(x���.[{�2#��;kb� ��������!�~w��.� ##����>��%
����o)�Aw��)sx�_BL�edZp���>X�K�Z�a�Ί��G��F*))�n0}�f0�#S���fp)����^^��g^���O�?���>����_�7у�dʝ�Gqu���B��G����c�P��d>䄃ůt��Z��)*��n7#�Շ���Ǉ^L�P��/� �k���p3u�3�eK��%T���P&��ju���"�n"}��Z��J�m�IwxG�?����`�jܸ�-���pՀH0�2o�Y J�+ꏟ�S7�����U��ߥ��2}pX����Ϳg�D�N�og�t��3-�0�&�
��7��՚�&<Q������b7���E��>>�/C�	 "Q�	0A� ���������>n���y��v�s�*��QX�\��c�3��w�H6Ġa�병���=�I�����S��@_�<�|�a��D�(_f�I:�!�&���*�d(���ʞ�e���fA� �&��|��Ȳ~������a��/�% ��?>~�[��h�Ώ�Q�FYz<���F1H�؅���������9˥s�9њ>�w���8Z�Y��ϔ��i�(Z7�y�˔1>�w!#�ϛښYFyZ2��� ɔq��}^�8�JR�J�j�u�˺�d5����2]pNc��A�0�����5���>���~q�|�Z�DlJ��͛����\��_M>y�v�x�|e��-5Q��F�wA 8e���F��d��r�?�0[�3 �7/7w��s�Ոs/_�쇜�Cv��Y(b��L�}�l�+H��?F��l��G<�!��ɔ����!����N�.U�xΫ?"ՠ=�W�u9�Z���G�n:y���J�Mf���+��R�"J���(k|�|�Ǎ`$�[���ܴ&���P��sr��5�̽�����6�-q������X˾w������.��:��<TW��r���/w
��}�c9�跩�?�=�4kT/[C�:-N9�Mb�^�:����NS=�̦r2�8�ߴ<\&�a]�~+3?��;.��յp���l�ۨ��G+//'�p�n��U�DG�ǡ�fl?��
 2@t;<�/O?���ގ��/�]/�~�^<��+�*no�=��X���:�ẵ(J1�r�}�-�H<�?₷��WC�ڤ�\ ��ۘ9@.��			ٯ��M��((�s��t�����(sd������ʴ��}�E?� �W[gl7G/��qD���i�f;?Ty�P=V`�PL,,S[�(sD���}�Jo<���$ߞd�a���!�_󾢒��[�+�p'�*|(���ů6��랯�8��y�O����V�6�g����zo��aK�pU�;Ez<@��^FB�^X�������T�u �����~�W��_��R��L�i����L'��'�"����8���It-���$����\^_�Q.m�0&�:�ڢ��l6�w�LoNV�fs��"p����	�y?��|��t>�tDĵy#�� TTF�C�~�=.�X�I������d��k����3 �;�����k��̾�0�y�ҧ��7�ԗ� ������/�;��r�F�Ɂ�f<E=�C<NV��>���[?��AH��ܦ��_T#Yb���q@]	#gq���OC���0�Mg0}.���a����h�L�M�j�]�0�K7g�o��h����;���r�tI���z��[α��q�&�X��2���7���rs�yZ������(����d^���m<��e�V������c4k41��!\o�1c�W�j�m"G��0�g�7��Չ6�9\�m��-��M��Ι��q��Wˁ�4E��hd�	Sa4h|盝��J�a���|�JJ}5?l��5u�����IN�`H�����v���g��1�}l�>g�/�R�K�$V��<���,�VVE���`����ó��G� �O���N�?�N���� �)%�U�m�\�dϟ���q��N�ct����.ׇ��1)py<��l}���ە9��F(����� ���tx/�G]�謍�(V7r��Ϧ��q�u�|͎�{gs��&K�?�1"+�d-}M�f� ��I���J���Z6&}r��y���;Uzϑn�h �����Z��1fc�� t��&!��F�R5FF���9r���H �K$���E�KZ�By=�m>A�[_�MWf#���4�`�����ZZ�-�!�rDZ�᠋���_��n��O,�w�#Fi���Y�G~FٸG�Z��Α�U{�*QW��s����|��0!u|:���9k�O�λ�k>;�8H���C��"���X�ɠr���@��G��UF��H�w�<~����-�{ ?�A�ժ�|�������BD��Ԁ��&��~���G%w�dɮ����tM�^1B�jmz���}�"C���B4^�\KyLIU�$b�͏-Y��?n��DP� �$b�ڢ?���V}�G�"�0Ԙ��i�5�l%-H[y�\�l�+�_/�~q�8nf����;�;"[󳰷������ǂ�+�7���O��S��X EJ7hz�<������	�y��tx�*S�" �*�����|�����N����#��m����a�߆ B�9M�{]�O��s��Ȱ1@�y)�k'�s`� �"ʎ"�9@�R `�h9Ef)��h4�5󶀚qui������0����7'C���l�7/�.%8
w�AV0�>���� {F5�Me�`^���q�$n^��_$3w��^_�|���ֽ�V{0h:��k��׆� G��ȿD�/�]��?���n|'##s��rS ��Un_BG'3���٢�ע���ӻu څ>���ހ�C�fcL` T��L?��ձ�Eő֖ cU���IL��4��m��T	�����4�&��� �VΥ'�����!�R�a�����7���FY�g�7nI��s��ŭu�:��s�Y�,���}�'.4��Q�v4ub��<�`��1�dT;QP-�a�{���i6����Bo*���]�~1F����ޣ�^�Q����|������ӎ���G�U�w�K:�����>�/���EccQ8B��[������r���oxS^��hu�3/77�,�O��J���<d�s�XNo�T�e@U�)��]�h2�t|7
�� "��:�[q��{��b�JU�J��AW�rS�3n%�x%�-�If�В���տ��S�N]���������<H��a"3OLP �mD �Y��9�D|/#-]��"FQ}�T����8���c��^]K��T�t��B�3�Ԫa��V��2OW>O�2���f��ټ?��bܧN|^������V��Ǐ8��	�����>��۝���Y�W�����}����nX����|<xuছ�1K��������O	���t������(�"S(�����QL{�y�L���#�T��ҿ��c<�9U��y�ϱ����re��ds]�P����S�Y��6�m�C���D[�W����u��4�k��i�8i����аg�&�[.B!n�A6�������v0��P��z��^�;�̞��m�]^]� ^�&�ǁ�8���t�qkz�-y6Df#|_��n�;K1�E��&o��WI� �1��dJ��>|-�ENɐc���Q����u���}�iDV��I���礭�;Q%V���x���I����Vv�������c"��2��o��x0{�6^��[�F�7�Bar�T��U����O�AȰO��������~d�b�--����R �Ah�I��@f���z5$b���r��,���E��(�3�HqpcEj"�oxg�T�y�$���UUo���T'��ɳ�PM��j3��d[;�T-�a!S�1�0R=t�"��$j�,��
�ɦf�"Z���\K�@I,��o����[B��%�B23�q�7|��+��������v{e�Є���N��w�h�2<i�e���>�U2��� Deա���s�z-M�g̙#�+~���#�z�1��ԋ������[���B���h���?�U�!�˲)I>�3W!l�pϓ�(5�v,V[�nQk+�o�����Q���>���,"qvd|r��1+R7���W�X3G��X����;���q>5�\Jm5H�R5;�D14&���P�|Z�����&�0�&�v;l�N5(>"`9�`�I��.�NƂ>`�&?��l�7��)a������61�F�ڐ��0��0���-�ii��pr����D�u�	_�泌�3ۘ��z�����
�Dg�5g2�~Go8����&F/��"�����!������#f����OML�],z��/���$(&�CaȂ�*	n����>t�ja��M�Q�e6@-i����`L��|3����y���q�m�8�4H�)c��!j8�F�<m��7�@%7��H�-�`���5ͼm4WH*M:q���!����֕�SH\ƞ8�L�t�7_=8j$����nK�$�0s���,�~;_ޯ�Z�5L  ���;sWmN�?��1x!��>p�H��͟�V3�!$�N��t�]nCk)eh8gnm�z ����l�yҩ{E���@�wb.�8Z�fM�3'�K'���=l�Lߑ��JY��[ϐ��5���*���/�
j��Z^�X�əS���7K� Bl���IDѻ�u�n��
��K�!fg�����?���RM��I����1�e�v��X���ɻ�r=���on�g��渣i�mpX��'̫�"�b!!���RE��o��Y�9�G���U��/c��eo��H�:'���%:�'e9O�!I�����Њ���ѱ �M���'7��h������哎�!AWL�sȴA�T=!��n����!�,�Ud�{%	#��Tz)	)7�h�$�mo�5�f])ႌk*M�_Ҵ�e��e��n\�K,��|I�1C�^�5�y��
�����_�G�uW�+��<�Y[{�.on>!��s>>�ɠV�tQ��g��~�wR�B��*F�?I&�A��6]��F�JC��c��fq�����H���n����r*򫟄ﴠ }��{��}��%z�O�Bߊ���9��7�r�����"���@�#��#+U��)X������G~tB��۾��813}-�D�,����7A��N����U�'}癧�ǽsu��)a?� �������ǽ��^^�����윜�:vcҧ�'U��/���^�ٸ6�#��Zr.ߜ�H�sTBp��f�l� l���+ר��S#���k���:���2���,<_��{X&Ơ᏾�R�$�8�$5&a2Uz[�n!Ǡ�����j^��)� �C�>k�
%�ݾ��Rå�t3H�7F��k��c�íz�^�k�ۏ�Ŝ����m��&�u=ࡾ���T���'B���9��`��VB�7���+ˉU�6@�Q� ���=���7��
o3�Z������n�����X,~\p?hd�rP!1����,�\��eސ�pQn�5%�Wi��4����s�X摨v�_Ւ3iZ*�se��������Z})�~���қ�����S��k�}	b�an�P`���X���rt:�ep	{Yr��X��ͼ�&#��mw����O�f���F�აG�g1p/��,�?~��0?z�Ҍ�\Y�ci��K%c^Ҝ����F�tUNx)�����
*�dz�m��C]�d�ō�Bh�z����`]x�<��������	-�p������m��H}�3D'��X	+}i��d؇K�zɉ���὞I����`��n}��x�۹
���o�u�B�5�~��نb���tI����霻@� Dd�i2��/l�*��L��
Ƣ;aC`0�q�Wa~�j���7X))E�����W��BٿN�Ԙ����XJ�A��ÊjF��{�\�y:h�_��%I������e' S�Kp�6�&{���0���	��SZ8��/PJߕ^��\5�[ڸ@)�>�$K��o��~��(�=4�͢�wYρ�U\ErU-�1-;C�=0j?On��7���c��;���}�ҶY��BAЗy�䆄�����A�]��r���Gf���!��*�Ջ�\���(�.6������Z����[okD7rK4�����WK�AX,O�&��K� �*V��ldO(}�ER����0��½�{Щ���Y+�&z��Un�te�Z;�C����U����PeK�{5�čZЊK�+���܄���y�/Ʒ�,
�
D���C2S�02XHc���R��u��9o�E��:n�k�v_R�h��J䲃5T�3�V'�ͼ����$�ʎ�Yq�>B����A��_SF�)�rV,llӧ�������Q_1H��U4i+���nlҧ��;�#��c��c�
�J�$��^����hE�N�Guh��H����1J1(����u�3{7���WN�;��߄4�0(������vT;^��O"%V�׵�U�SG���tդr]��2W��{gV�;��g��n��*�%��A',P�r�	W|�����&3:]'u�� S��&�=��fz	��6Gon���D�U��:~�t1X8==}�l\:�w�Pl���A���b�	��V��٪�:ez���e�|`v���.�d��%+b�<l�|V�'�廬��d(�9,����v,�s�(�fm�=�Z����O�,=��i"�$��@*Q\'����PI���gMwU����239���O]	�o����U�m��kmU(��ʗ�#�l��$/�{��(�r##R��!���рo���E���K0X$GőѦ1��j��mɔ'��i8�~�����v��� <v}s�P%+�����d�Z�,l���]�Hi��������k��������Fb7�%���[�O�#�Js��*��:�l��b�4�n�eݔ�&)�h�s=/Վk�,�l�r�W<���+u�\%7oh{����L|����UJ�2���9�t��%�������\X�d��V�'ޓ���8�}��섯䋘���D����j�pO�<"��'�_b�� >y�����P��g�s����Ƌz���&�1�\j/Vl}6�|��� �*OdU�K�����^�һ9�^�����L������k���I�2��N�Xb`cJ��W�\�C��SR)��<�:w����M�61��4o��Gއ��p�(������}`7�����qM��r���o	+���U��;\ҟ��׺|\v�S�߬8߬V(�����r"���֒+�'RHx���)�U�	��=����E��l(�I�/��94��Ȑ�NPks]��rdlgg�t�|3�[tR�M�"G��Y��5+5�w��y��_|��,+��h�v3'�&{�]�8��^`��6f7���S��T�f�Iv|�"0?D�B��f��K�\_�DS��,H�U��W�=N�lڅ�>����~��YA>�O8A��z�XA��vC�#���{�*2p�p#C�Ed���������w b�XæF�����ʍ5�B���P�{(�	�K.�#�nX�;��$=�W5���iF�>h�O��	\�(_�nB��[u�c G����iT�*�����?��2����-��;w� E�;�����nŋ;www�Sܽ�w��3�L�%3���9��n6~6F��6�5�͐R��~o�'ǗZxh�,0`��������>�?tl����I�{�v'z^i��-�~*�����5}cegj��w�t��?*���1A�Ű�83�m�'w��I#�ad1a�ы5��5~w��]�߽�a�6I>�s%铃Д$���3�~����2�.Ȭ�jɤ2�;��$�I�6��DA>n>;���Ӵ��vˆ�wIq�����Z�C�>����j�N�����AT�̼��*<�0�`.���6���;>$��q��_P�9�Ȣm��ͭ�7n����\���ש��5��w�+ɚ�	DM��-�i%f�Xq4�W�_>q��%H�������N�6��0z ٯz��|�0]�CȘ~��۞?��c���� �+��)N��'����qY?���s�̲��|8�
��O���F��m���/�������n�N8��P���3�~�nFh2�v2�ʂ/����N�D�+&^��R�|ݖ	<��T�+�n&)�j��:�EM�<ƱH�<�����Z��c�k���T?׭��MX���i��̭g��-���bVLL̝���V�EyE5��G�V[�Θ����eG�mI?7�<p��m/�я?��8���� �>�L� g>�~V�?�����j,0�$Q���b��ᮊ&D�2�ڏ�ܷ|�YZ/ ]���?}���b#�{h��ˑ���N���������"�+�l��?��T"�y(��O\,f1����̈́�:���
aɗ�'�O�Y9-i�fѦ��&K���DCz���"fU�:��f��ܞ�����K;F�ьZ�L�Ҝ�բ�G����@�Yw�s�>�jJ�}+g�[�	����$��B1�|��$�5��7Ǝ|u:�]�j1f�j����y���.m2�)�>Q~�"F�%ݎ�p���OO���͕�lB'&<Tht�^4�oZ�B�_N���M_~r^^$Y(�t�tQ-4��#�<��`���^]N 5�5�}(}�I�E�ՂAt�JN��׊bZ�'v���*4��C����4}
>�xTU`���*��ւQ�PZ�k�V�S[�l�?X͈w���c�����;���10,=�N�2%_�#CYUʘ
�2(��<T���g6��c�R���M�s�0���w����ZUa��if�{�ggg�1x(��6��!I���E��Lģ&'�{Wxudk�UkU�޺��̒W��n��n|5��[6C�zTkc�\����݊m:�:�1w�%��ׄ�p�k)�J-�:��9��m�V��(�֢�'�8�?먛
"��������^��]��=��������ml�'5c-/Ӫk~wI���ԇ%��ƨ(q�'�ᱹ�=��l��O��'�H]HG���o}��V�T���M�.��p+�M}�n�A����W27*���5Uh�X�I/�Wi��=B���B����+d��2F}ʍ�O� .ҬA�f�[T|�]N��ML͋X����+����>����<�t���;�'VzOnK"�q 7�@��(�]��i�A�Π������'K���AN5I�;)�^�7�7���0'W�L����pI�6zO�	} Շ�I�VE}��T�q��w�{�e9)LwA�`u�L�P����б5�1͟H�/������32A)��d_��CW�dd/�OK��-QW���Yq�7O4K�?'�۾���wA�W��L#.����� !�^y����Q�쇸�Z���f�g>Z	�r�(åD�*m��m�Vz@H��a�&Ufj�gc�$�?�c3l7���E�mPK����pޱ10JH��Q���R�C��sΡI/4v�U�Y�@8��z�Ψ�����>v�GD7�9�S�b�V�3����EDt�e�+$��BA6����WJfPw�ŝ�q�79pT� �d�^��V���̖76����Γ��D��H� <axs���""��.h4�M�`� T����ϻV<���4y�YN���t�׋bOJq ��+�p�~M�*V����+�^ӺG#|�uP�ZVVó�70�G��㐦LPvXe!=$��xq/�z)a]=����m��EI?x	��RC�F��C�E؜m������ؼG)x'�v[���$������ɵ���TʘiJ��X��+��d/�l6�t�Ro���ΜWD�T� ��T_;,Bn���v���G��fȍiƮ	����q��b�o(�ڌD�'�v�1�&�8]~UY'sr*�V�ԺU,�wsO�����s+��G����F���֡K#+g= ��8g���X.�/͔0X���v�~%)J���b	�YH�S�D��B�	��L~�V�<�b��0ɟ����]�.L~�A����*R��#�Bq�Ԁ�к�3&�b�P�Ee�0r_�y���������o�"U�j��'#�YF�K:S��:E5�1$��e5����4���͌Q��,��9�����5�&�9��ť���w�	ܖ��D�S|`�[�i�^`���{��ʋ�ZY�բ�"�s~��s�A5��By�ߗ����[2lȠ�MI�K>��9���<���X�D��U|�����J�ƿf����&��*Z.��?W�4�T�!�PEz��n|���ŐG|Vy�@�&}M\	����W�K]	ھ��Y��!��0Ox)����S�d�r��/�KKO�4ag��8FAH�\�I��>=hsu�PK�������|��e�S@��Z����;[%�}�U	ބ<	Jn��0��B	����f�n&�;�vd&FT1oE�e������_i�*���l�-�����l�=�[��ַ���Da3�mfw[�hu��"e@�V�ş������P$��M����ҽ�M)t��ɳ��Q��S���) �h�j?s���ױa�Cx�+�bb�Pv�!2�o��b�4�;SH��(��\ ������W+������8���885�������)/�v�x�����PpcH�1*q�M�Q�*C��JV���1�A�2j ����碉�o�仼5hd+��k豟sc-e�[����~~A�<�Ċ��:]��8��e�%:s�4����+������6d�e�f>E��u��[qk);�pm��x�6
x>-g�4{z�4"�s	���|��(��
a|�f��H0�W�����{�,�� �x;:�ggg)W�����LOO�	��e�r�ГJ~>~I����,�锚�Q(2@��s�"�V�6��z�%[<��9��>N��P�RZrRX���
�L�7���2Lǻ�d�|�*\�?nOY�a�I}ϑ	*K�k��V��ϔ�+�a@(�pY �`�M�d�CN������Y��XY?�s!�߲�2N	SX<��"e\hJ�������b�֨�}�����sX(%c*i�����L�M�i4 IСHOɫ/LL�>@.c��D��!ڸow��e̬&��L����-�ǅ�H��}�e�m�͌#8�?��d���H G��
���	z+$߳�zy�#6K�=���3�v��$vvv��sGYk�����ٞO�4o(Ұi�g;����p�:�l-U�Jb�^����"�(�siBq�%�<
^�n��r�l�N�Z�$�e��t����j���<ȅ�-����.���,�!:\���9����(�o�p���*����ꗚ3����\�$s�/Nu]��d��\/!n��o�/	KW�i@2e��)�x��EmG�x�h8�X/Rh����I̤D��u ~+�O�H��0��t�/��W�4aQk�O����H�5��]��β̠x��3�!�����@�U��^
���Z&��f��I����0_#P���������	tOM繲�~VF�/��H���Ł��V1�T㇅�D�e�>�V��-JԚ���z���T�k֮�8]��͑}e0XS��F�����س��\6�~�Mx�Z%ڤU�N����6ď��T�ē���Rݼ~�q2�C#�:SDh$���l��A���[��ݩ����`�r��3rӠfD:Rq��.8`!�g�r�r5�=&�U�[$c,x��},���L���\�AA$�^�Y�뗑�\�kĊ�?��O��?�vGHfu���<�z�Y�w�>�������D!{w"��3��]�#U��`� c5~�ȁ-d1���܄4�������k���4�{��5�{xn�Fi}KW�G�.�LB�|����O�����>e�	{��MQ�Φ�ҩ����ܘ���'�Ёr����������}K�䜢Ф�_���ЎL�4�hw�`T��S����8FZ4>&^�ɹ�*Q����{8����v��*�*y5
9PX��I�,���L.�]��A�'A�\��B�g|c�0^%s�����S;��F��K���e�"�\�+�D>�Y�&�1؎��ʇ�Wڗ�?��ie��>�M%y���	�������Oeu���h�6��-�X����&ֽ3��|�>��# -��ypԈ��d�������8^��/��駬� bTC5d,���V*؉��{vYr�!T���P��J��x��=�0��Q��h-����R���`ٕ��p��e��'��m�W�=龍|n!a�����wf�N��FyQ�����B�H����#����X�v;��4rL�s���N"�q#4=S ��zj�"WO���ki���3�M?����ܝ��aM��>
'��D�ј���a������X��?�ʒO��Z2��<�D��FiմRs��O��Ef���,�OQ����>�BSE��ס:r�pd*.&p�̲%X0��΅�Ӊ�T��6>��gH�J��y�'����Yb��R�%|������!�;Ӯ�юfûg��%J�H|[�G-"Aِ�0>T0%����Ȱ����8����CAD���w8Oն��=&F�U-�����τ	�?�K��UW�i�>Bg_ۨo�k�a�
qy�;�	b˷���ST��"�fĕ��r-��vN;c�_r�{yB�.�.h����q���d�k+#��R"~9Jǰ;Z58�
���Y����f��ڀ>��&�M������|����,�c���a�9�nWE2��K���$�K�����e)�;���TF���,E��7�v�h	����{q�E���nإv٥�9HUC�vQav~�o��o���5K7�*^����!�W=�����4��#�Z�'���|�(�e�3�,X�5�&��9��p�X�G�;o`��6'�^�O�6if,��4ØOe��i��!|P��s�V?+��
7���B[�v�W��i���<�T�@����>��:!PF��=��i�k�2w��R^����V!���O�VY�s�������.�PL�gEs�h�tw^��ٶg@|ˌN�(��K����dϋ��ǁ���%�W�t������:�._��(Fqs}?w�[g�^H&f�O�[����5��%���%
���ar
�Ŭ ���g�V�3���R��"ٱqp4S �7X"�f鷯��w[��U��|8?A�[������.G]h9��E��7���c��{��^� �X�0 'Q��$���rk��[X$ٿ.�qvx(!�V�~g A]mm�����F����}�m�(C��Ԅ�ѣR�N�X�Nk�C��uB����P��p*���X�@��R��g��"[�-�����>f�B�g3i�-lUKxal�.歝�T����@�7��z��;_�I��Gq�X��S�e,��۷h�^'���,,��#ۦ,VE�_���x�ͮ�F�Bi�������
�'	� %{6�g3�%f'�;�����k�XkC�1T��O T����{==$�%a��F�_�z��]�j��LԦ3Y�	�I�%ʖM�|����޿��W�8���Ic��-K���V��Ϲ����7d4�Q?��fg����z��B�I1p>@���l��r����̖h�����˶��2��3!������w���_�η7�H��kM%�6t	��@"�W��M��Ժ�ʖ����K�n�����
���t�,	�\-}�?��sICW��}��(3�sYo��:����&
�Y5Z)�a1q5��*g�J�,)ٮ㻳dHZYx:��U��xC<Os\�Nv�/[m;P=7|=�����e���w�/�~~9�~3`5psK�����Tf��v"�쩾��!O"��2k��]��(о`��N@�b���������y�#�^���NJc�ؘX��cƒ��R��Kn�9�HhP{{{S���^A���u4��6�W����E��5,]�m��|㾤��dV?+�-��.��/Hz4AJj8�Aᡮ�I�ӯj�P������`]~'��͊d˫����s���֯�,oŖ������I*w���jc(�YߝÜ���j�}jʭ������:`��n^��oR-#�ҁ)h��j=W蹴ç�C��κ�ԇS������<��X;<,:_�c��M��څ����\VT�U�ަ*Td���fU����Rs���.��^z#�2���I7�,�Fs���0�ѩ�u&x��e���@�7=��K�\���PD\M�QYW�މ	9A��/��q=�����|����@�a�06>>�O��	��L	6��5�ft<i4�%+�t�WZJar�D����/�.�Ӏ]��a�x,��R�KR1������dvD9��{�{�b7PK|ފS���<*�&��?%}�+�nys%�2�,�(�a,z .��[���.���-q�T��8�����쁍(�U��#�Dt4���/��-V�6�-�Sf� �R�ת�(�h��yY	I�C̯d͖l[�wߐ�}U@+X ��h	FDF��{7�ws���+���鬝���[o�����?Bg����CG�|kɽgXU�٧o�V��˒���j�����2q�c�.��ոȞ�ē6�~L82 �=������,,�{�C��mr��F)Q�=8i:���@�i�`��N�[��^qBdPN�9�b��Қ��_��.o����<�
s`��t���ʕ�FZ��QY��!��y\m�;Q�!:Ȥ�Z:v����<Wb����~��笋�=n�)2�)����xl<_E��K]tj��YA�H(�V���G)�,�LQA`ˇ��R��í.Ǿ.��*$�]O��0\��*6��ۨ���*{��yif��_�F��Z?�=����B�����)�Ｒ�F��"�h�{D� >�C&�r�]�����%,'�P��f��� VnS+:Ş=ňˬ�}t5�YP������������e�<^���#�h�����+��d�?��M2EF�I��s��C~|�zD�e�"���L���wN��&@f�m`MnLf.7�W,�o���Վ���������F��~b��)%t�*l��'��U�0����0�Vt[���ew1����%J���M�0:]�}g����7Eab��hƙ�J4sN�QL:S��ʔ���}�����;���F����r�'�~g,:�5����"�V�1I�q��)�kң��Hǈ�@,����T�9���I��e2������rǽJf�X{Y� �h|'Y<`z&	EB���.ϿE#<��y{G`��M;�e�����}u$=����^�ނ�����Hk�/Ɖ��Y��f\(-�)�HB��hvw_��عU���<�ؤV ttps�n����z��s�8���ƭ�D�l���nuuӫ��'+U�C��V�D�ПN$UjQ�77��|[Q��l���2�y/3�8{�zz�¢^�g�j��a>����4��F4- ��W�6iU]�E�Zw�6���i�A�<��KI�ڰ7`.�PE�Y*jiI4����� R�A����sv8��w��$����pc���NoY����%�)�w@��Cȳ*��S��;��4�9*٦�w���a�� �296���l�����/���g�E4<(C����}^�V>����M?H$��/���]�gx��zV�z{�np��[N,��-ZNMV����L/���2{��X�����o����z�ۚZ��/9���W琧�X����sE3Je��$Hr��:2j��Va� Vt���z�'-6�R�F}� `S~� W�5�0������c�g��s���r�~tq�F���8��X�e�>���b5���]�PNY�I����F��NO����|�����#����X��`G�����p|z��g�P��O��K��,�,��+�~8�����+��ΝoW��.�x��JԮ����$rp$R�ZU��:QCO���&3�8O�b���*��m2��<qpy]��,��!�l˙�LCC����t	�%�����Vy�ݟ弌LL���?��G��	��wh<��G�qYu�!1�"K�7 �7����9(η�,*Q ܰR8c�f�l�
��_����8A�v�,Vtl�Ř��d�a��Y�o)Ɖ#Io������ 
�zd�oT@Ѯ�@֛T��ʜ!R�>V[�q28c���}�T��@��'�?�j�ff�H��K�^��'Uj�4�UUeLȎc8���t��~�3�h��'����B���0���g'i�R�oJiӌ͔T�T�	�X��(ƕ����Y��6-G��*2���-�h;2�#����.��&!�2�^\���=��{�����j�	3�HSn���<7�%�:�uZ��ύ�P��B{oDC�Y[Z�:8�vZ'\yU�9	&��de�� ������ʜ�Vd�`F�ci,#M�(-e×�#l3Ŕ~l�I�&���G�}G�gJ3�˭�Xg��]=d�v�ғ�e�T��tT�!�ML+3�B�"�`F��v�Uwqi�fz;Fo�*3;[\fԄ���-vEq����-ަE4w�_;��L�� �sbr�HVx�io%q&d��By���a 7��|`4�A�VO� =;�<U]7ܯG�]�SjkcC���T�b6�b���E �v�-�;ᚺ����,����($��-��,=��
����-k��,]�CQ��Mkm~5⢴��*�����p�i�A�s%�q �����$����;R�i��E�Y�VS$x60)n���d�`�;��{s}��{?=*��b
]>|$�8m���l/��-}��x��W��wl�/..��Y���D��#�U=�gi��Y�`��,��}��o�xa������`#G����:\��gd)�*���.��*.I5PG���7s�GV��G����� }!�)uL�����;�U����H����X}���Ł��=^����Bne����������9�u�uLB:6�ē��
�B�[���&|6���Z�6׈��R�P]��w�֩�]�%9O��~���4�g�j��®%����BSs( �~�*+x�Wed��s�֕�!�5�	@+W�t#D��?�͇n�=�{]!�����ߥ�B��B7�/B�Q�B6���'Ζ��x�d��H͖�ײ� �8U<Z*k�p�z�_ �.�Įl�|R���7X��m.w�4��8L�m�����nt��ݑ�ib�AIA�%
{qa�jjjx(�|nѩ�O0)�u���1�@�ؽÛ�
ܧ�D�@��P�?��|0m~P�y��;>;���H�4�����>DQ��޶>�I޷�^�1����]�r�������_��ƀOT�n�f� �*P�"��Xm��a��PQ|FڐrnW�����͋ڏW��#��읺Op�������_+���{�k;E�)�N�s�<��f��"�<&�sd�,Hk�<vO/T��$�(�򠜞�����y��2H�ea40�]7��	�r�)"�����"C����?̐�oI"��H��X����N�kQ����,o||\�B�\s��O{�Mv���u���4<�����GՂI��������K��Q8��[z ����B� ��7��׷-����s[�ic33j�20�8�w�w��Xq{��L��<c`pޒ�3�1�0@>��{��=W�����0ͦ/���߶.������o��E���z���<S�,�h9�8n�n�n2��c�O�+q�[��R�Z�B�S�9�BQ�v���T��e�.Ԝ�?O��z�#��F�^7�u`k���Z���U7����j�����,�!=;{�N��gz�nGeކ]}#`��:5b�Hljkc������5��|j���z��cy��(<ׯͽ*�������_��`����z�G����.�F����șs'��'Z�n�KͰcE�'H�W7tv��>��x]�0#��*~L(*P'�O}����v�%��Cb�����1v���`���j�+#��Q�~��&<�t��*�G�V�� S������Bܦt���Y�܃P��,Y�My��@��ŭL��@`���9��fۃ���^X?1� M���	�b�aqc92�߿��O�o`��QcCO��0���>�����-����R��h���������'&��>����\*��B������ǲ�o�o�F�����H�1=��MG���Y����A^]�{t�c���7���S�䊝������/��ۜ���Z�W�y��w��E�N���x�e�ic!EG�!����vz���/�Hk�AW�m�=E"\�P�����q�D��]�������?=�_/�\��a#|8V{]�ߧ�/����)�z�%��F��v��E�g���9sq'�縹�o���_�������9uey���9�2���qin:W���0�I���ˈ�ʩ! ZX�g�_����pY�� `bݪ���n�����}k�S4�8��5�6�C�X�ؼ�t�� ȐT��:���{�9#��T�9����Y�(5�)�]T�$��	����a������9XǨf��/o��'�����p�����)��"�����ҳ��xM�K8;?G"��!����Ifq�9��B"(�4�����WbD(z��P�`����%L��m�l��P�Y�S����f���`��[!o����$�{.@髻���`=;��� �VEk��vF�Ix�u�(����\[䌅X�M$y�N�u��S����z��嗶3/<��eHbX�\��U}�;]����Vw���Q9�454L|}���S)c�&��[���m2����;�ӛ��j�ܭ.�|:=�17�Ij)+]�X��y2������:f�-�F�.�5Tl�$�/� d#�aT��a���n��>��Q<z��"��S����KTD1����x;p��q�X���`�}�Ǯd��1F��/����3
!#I �/s�X?:��K��l�"����]�|��n_����+ǭ�B���d*"�]u:
�ֶ{q����4�����,�9�u�XŇ�II'��D�K����	����=�u^M;�g�\ߒ�r����=N�N;�7�;��V�^ɲ��J{J����`��'�||GǙ�j���J]�l|V�bKQb�r����`A/oI/��u��9Wh\�}�cĠ4)�j��C8W�Fo,-l����^}����u������y6�\�ް;�_p'2W��o���R��3��F�2���S�Ý.���l`j�u��O�����a��N�9�����?�P�P�6�0l�1���1X��>�?0k��2Ŗ-��,e���0U�U�hi�n=]�ۤ8�ʚIcK�֖�A�p/w�J�A��y�m��c�>���@�$׾Lābɿ��;�*�*���HH���_�/�jz�s���{�6/p�}�5����GkÍ3���t�N��F{��>Htۜ��@q/�������[�^?���<]��vݠ�c67cYO�F�T�z�-�0�L��%��:CP?�r����,��U5�������sm�s�"���B�����@>c��v0l<�H�,�nU%�Q�m�CXN;Tf"/���a��U�2�(�KFU�]C�bL��v%0L�i�|�+�
m6<^�]��4=g��u�j�D�����7���*hOM�\���-IlͲn`g8���r��p�@(�8��s����<�*[>��/,�S��䘅�{�����=�E�=-	x�}�������(�,�U	�by�g�%�b憡��Щ��
$]�1Ԡ�����rI^�@BO���#,�o�qY_ �:��]1�%���}��V]���/��1h�D�h ���92\�g\#����ttb�"Uす�gUL2S�>�`���44*�>�k>hˀ@�_*�3˙?�����Y�U���׶��..P0�("���:�^�eY� �d/J8��G�Yn�W"OOO7����?�m~�#y&���e`-Yl��"�e�J�@0%ˆ륖
^}�y�W��L������������3���������\���ja��-�V����p#I�T�t��'���G���~�W������8��e��K�O!��}2Q$��y
ټC�f��Qv-QhAmm_WϹ ~����l���xB���PY�U�����!_-K�M���O��b_��P���.b���C�\�zJ��{<Q�4,��×*�j�rwr��lk5I���l�&���hn^�T!� E�%kh �?`;�9���1H��*'(L,-#&�u�.%��)婒eB����^�5;�b=������:f��++�h6u���bq��u��q�x]�����s�wGw^����{�lC����T��Gqa:>o�~I [���[���p�6���%4�+$���=va���:s���!���"!h��m,�@�8�'?���N��z\��b�m�#O�O��;#�D�� �%� ^a�`"X�z�Ћx삳����7O�����:�B���_c;ÔQ���k��٬b{w�%����NCj����g�Xi��>����a�;�̡!qh���^���'w� �C>s��h�Y���`Y�ܳ��eE����))�x�ϐ��t��Ƭ�]��a�.�B��ߍoX��;I#����������&Iҡ��қ�.�։��j�*���S�g�Vo�Aw��Cx�Dx��Q�=�ŒZ��9�z�O���}�f����ܩ�tu*�x(ԎY	2�����!�"�pa,1�39:��
�v��͍��D!�B�������$��Ѝ����ښ�
�Eb��d������$Yф%1����@	��:]a�u���5��Yiv���3�6E$/�b��/3#�kK(o'+�)[�Y�#s�1qu�/r�D���]���dFw�s�m��Eۮ�(�(
�gͥ[����c�u����nF�bҐ��F̥�Ʒe�o2��"Z"�e�.�58�֛�LN ���њ9{�o�"?Sҥ�9ت*����åk��$���s㡤k�n��5�h�~`�4�E�'��΂�N\�C�7}��e۰2�j;/d�Mu��[��ѩ����C��a��l&<�o�nq8�Q��R��rm�x:{4T�8�.�w�u·,>#������O�sg��|�|��6{S�z���W!�̨��QH[�N��ZЮY��9%�/�}c��N��\��eL	q��ڤ��sL��/F%7&�9�#U����s�0�Kp���<��~��c}�7߻J{z�ș�0&��>�пg���P�M%o	\��_�a)�Q^Z�[�xt��`��9�+���y�j冟~FW��T��������Č^g�Yx �`OV�BVT����|� �Qc1�j�2E.G�ڽ�D�ݑ�eW+C=�u`�7OlYJ���m�\"y� �\�qOOZ�Zy4���X�V���q.��������&'J��bݥ�˝�r�$�H��a���W�h�q����}�5Ѫ;5��D`v�-�(�9S�,ҋD����8md���94a:cL5k�v#hr���	�lY�(z����$�X��zJ�}kl�mY۱FgQrRxC'�i�j�}�k�7�#1}X�-k[���$����S?����8m�c�P쳖�/�rE�hE�z0�`Qΐe�T �jq��bbu����S�pn1�y��es����ï���,��6��l�4�u�±޹<���k�	�<�"��(�8������7s ������(���,�B:�Z�V��8��ā;��/
g]�\�	�=�Z�nT���9ު��3��2E��XQ����
S]���ܨ�sP=���`�2�����Fw�!�h�6�Ro�su��4 +��cw�V��WWG��:Gc�ː�t ���˛��	���?2�n��k�ٶy$�g.����^B�F�T,�I ���6�����+Q ��G��(���odn%�Ⱥw;&�c�S�����˥�!�wq߲�t@V2���-�9�h�3���3��`nY�g�wy����m��$]��wN��X�b�_���/�-1p5�#3�8��mw�PӒ?%ٿڍ�!V$�,)��iAͩ�FW���X��	��g���r�(�"1�tvO�4�N�sH��Z�2&�bY�Ml�\p��8�A�w�>�o� *�I�"�8�_M�#������&<�����>S&�4��'������ݹ\^dbno%�!h����� 7�#]�W�L��a��P�pH��0��\�d�m[_'���Z����i�ZH�[91""�O��B' ��gA��O�=���Z�/�L�t�q�xH�������E+��j[%:��gn=�(�Z�T�Um*��:z�p��8�cpH�m�ĀY���/ұq!|]�n�T�u:c�~�(�4��1I��{�o�b"f^=�lEbH�U�7�����"�nk� �tj,P�W�x�+�������D�(U�
i���9x�q_&=&�U���j��+�p��ɅM�i��!��LW�Ѡ�N��])���f�e�@�7�І!Idp_�L'
���1�W^o��Yy��e�m���?��>j����ESR�$����Exu�,�pf���^X321]-�t'0�|��!�q̝W��9o#X���g��w�NNƖ�S�s�s����_��E��4�+�� � F��8YU�ZSS�b��Udʟ�!p'�	��B���jtk�liפ�3Y�a)��Q�ȑ���)���l�P�e#�s|1ݥv�|(���pd˭��C�ף4e)c�����jz�������ݽ��{	���2[?	����)rw��ާ ��q�%�.�ŞcCگ��R�z5�Uj��#S�u��΁Uj�MZ�#R�������\�ǡ)OO�!@G�eu^6����P>.�"��
-����R^��_��* ��h�v&��N�3�r���ڍ����{�C��^�<�k���p���2ؕ��~D4I{J�� )��aL�V�}'G���#���O�05��6����c���Q�ϙx{g�U��ࠚ[Z�� D�K�I\-Z�_�Ga���
)��"8��.\w�{"5���!R��_�6����ҭw=�N:�'=8�F���}�����\����'������	������s��D�P�SR*XQ"K�;����.�+�y�T������E�UO}����[�����[�[�O�?�
�M���d�R� T	y�+�8�j6�-�^��j�CT�H(7�������Po\��f>��[of�GBL��Mră7�.��sR�u=Wi���	�K'�Q���C�%��Yh�����,��w('���~���r���EɧO����(32�V�
]o�J6��{� ��Um�����?f���]���nұ!vTSB���P�^���s\�����}�p�"�>ܾ���m����@�g��>��P_����=V�'w�M���7���lK�X�ؙ��J?�f5��.�m�2n`�͐r���89���DK�պN�ء����~{�BOe���k���u�9d��cn��%�㖍g[�9��49�ȿKK񃻻�QQQ廤�=5~�C}��Y!Rr�h���3V�[��͎k���${^݀�Rp����([52Q�j���?T-X[��w�,�"��=���dEZ\\���0��K�i1�����I���>�Wۢ����0U�D�j3!�3�>e�l<�B%W�v�~	�D\>��ַ��Z�JϪk�@Ғ[G�i{��⒝���ԖG�Z����W��(7QK‾q�
�ȡW�.=k����QN��ƞ�Ƿ2��g&1�w�ѯX� ��:O�w
���	qފ
x�l�
Ƞz���^d�;�U��r��R�{���Ln���};����tz�j��wf3=w9}� [:;'655eEc��gffBD"�@���8�(�Ѹ\64�UЋ��ަn��u��_8_4觋�=�;�C� $HL+&P�{�KJ������6�,t���}%�#a#��\��i��@�G�����U�5��V�;���'�/��1�F��O���0~�u�]�-@�!C��M�A��=7�AUĎ���&$���H�DH��%��EJu�'E���hm��� b��n��\g�r!��2B�6��b�J%�H�X%�X�Y/iUlE1I����(�qm�A�O�\�3�b4��nUpݔ�GzؖK����� b�2 z�i����^�i�$QJ�.A�R�*��Lc���qf�[�F�j�Q�TH�A�n�U�c�C����	���)�0��P`:u���t�v	i����b�R�E�Ӓf����}X�����4�X�*JlW�.�0-��d�_d}}����#�x�	}�Qj��-g��%��o�[���C����2t��^-ځ�ǃ�-��D��4M\�ʄ	�]�ڨPkT�T���Iӈ��1�� {_��:��"M�:��R������v��=3�b4��	���rU�@��#��h��y��@;Ƕm�l��q1	T*ayyY�.ʀ��OS\ۄ�v���'
#�E�eI�0���׫���T*Ah��s�q0��!���:����B}�h�PVȃ�����l�a`����^����ԛ�\�pnFQ?����o��?����q��M;sĉ$#l�D�*ި�.j5����dr���o|���2á��Yaw�F�R�Zj`U��kgwHeH�^%
�*��j���ʏR^� ����T*�!X*[�u���������n �R)���O���[���`yyY	(���.+++DQDw�W�7)%�dk�:�e�x'1�SƮ9XV��q��0���E�\�U�LS����U$�{��#�u��Ϲ諸U�o��G�D�E�E���3�ʱ�1��$���$�^ل&�&�"@6Y8�d0�ăh�I&�c�2,�{L�"m��~UU��>O�ۗ4�T]�
� |4ϭ��s����}F֓�#Z->�+��e�֤���zY��EI��k�Z�^��0�p]�;w�G?�	��/}�K�~�"wn�&�)�i�c�ʏ�7=B�R�0(�H�L#k�?B&�c	���7�Z	��m֏��?�c,L��0A�HbI��yP�F��D�S��K鯞8A�QG�U�ya�4}�q.��aN�(��u�I�w�!�t����ȉ�8�J�G���p���40=H5A���[�6#)�	�j�1�ZI���z]ͤ2��޻Gݟ��H�n"�4U�2ɖnt/F)RJD����f*���x<ƭV�Tk���U.5�ط�!��O��.}�W?����q��]�F*��G`�T*�Iİ��^�id��\?WG!�n��O�������'>�������m���$XB>�U��	`96q�0�#66_�0>��#����kTj5Z��X�	P��.&�_������&.\��T�	'gΜ����� �kд1�uj����]\���5^z�%�߿��%�vU���l6����������ɣ�>*���0�a�!V���;C)C��+�A
��x����/�������	���p���u��Y�k �m�L%�h�1��0O���((�I�`}�{�GKV��y�3�4��#N�<�L-�j5���}~%���eBO�-􆋬�B@G����r��I����nﳶ����"��V^w�m[	Ogan11W���J�QC��2T����&v�S]~�g/�η��J�?%'��B2hu	{�c��wh��sok���e�c�� ���6�qH���N�����9���Z��NP�I3
���F˶��gϞe4�7�8?u�~]MRk�����P��y��wI��Sm#!��1
�DA��)�s'wn�18�2F׭�oY,/���ɂ����AL
� L�D���2Q�k?f��o1d��8��WU����*�7_ckg�ᨏ_�9~�87o��kIE�0}b��a��eZD���BR$/��"պ�aܼy��/�b�)�x�iC旚[��؂PJ���?��?�Fw�E}q1��JS���}��a� �a<�a�ק<<%�[���1���M���>�0J�Z��ܺu��}���0vk	�2��lp��\�r�o����B��;ɘ4M�Pi�����2���S�c�;V�IV�W�� R*��f�cǎ����o����eww����4�ƃ���vH#�(ngo�V�E��֔��:=V��4M� ȣ;=���\�É9!�c#b���_�9�u�V��a����2��I�6�iX�Q̉��p �6���t��F��82�	v���ؘ�E�WM�K�����gz��Q���̻ex!)�L0=��8h��dt�8Qw%��!z5�{w�x�w�8w��u�kN�P����y�p�{׮���!��2�0D&	�e���`��J1
9���� �˰iz>{w��̨�	�шz}� �#N?����.B*
�h4�G���cG�qC�a��!v�F�v��k��`���O���2Mj5���}<����$�%/.����-�����V�E�9�p<���3�;-^|���9�����C��0BP�}���XXX��HI!�j[T���R�$������Ǹw��/���w9~�,����I���p��9��ܾs��AhJ�~ �6��v�� ���H1<�B	��TeA
HD69]�}�fD� �b,�����W���A�94��*X��Ƶd�V�0��Fܹs��8�>��I��4�sz�Ƈ�oߧV���UfZ�R�!�l���Kc��G7>���$���l�ߺO(G���,L��a�)�r�������GW����]���uKU�ۭ��q�zD��iS��Y=��ضK�a2��K������������v�o��t9��
g_}����g+�z=�D��秋��&RT=�,�$�0T�F�������4���9d0���+�� &��D��	�_���[,--������I��n��1 ��K��,��F�US�!�>�i����:[�c���K���a���UH�'��,�y�j��e�� ���_�3�}H��� �0�"bէ+@�b`H�Ȕ�D!�4b�s���2?��x&���&�%	��1̔4U����/h�]n߹A��2�p�����$2&��B�����1�G�������.�N�I��ģ�������txU�URo���wh��BQ=�]����4���w�JBFq����I�ʢ�:�,�J�cm�8?��2Y�ۘ{�昛���'q�):`�)],�Cn��(���XY�N��ad�Wf���Tƪ�t��F�.����m3GHT�EA0���f����z������j��=��m`��,4�$��4I��$���H�È$N1��t8y�,���"���[�ܡ}0��X^�(6�1�tq�
�b���G]�$ �F��T��>�h4bgo)^9�*����%��N�K%$�Ķ�<l�!�$!����7	�1�q�51��Li�����dnn�n����6RʼH�����y9(�1a4D	�a�Ѩ�0b���[��s�c�YB�D�iILK�7n��f���-��:��~���$ID�D�1$���k�쑪�I�5���|R��xj�
X��EE=T���j�
�_�%<� RSҬU�l�A�mJ\��6!�c��׳�*��K��v��yY.����Q`�:s|�w�k�^f��݃��P`ul�Ǳ�Xf��iT�z��5�2����D%�eR�UU�!�ٕ�벾���ٗY\^�Дǜ�!����\u��J�e4��u{�j5�{�.��ַ�F�͸B ����8�1�(P�L�ƶܼ`x��/�T]N��b�)q2fo�>�/�´���R�T��eY�|�q�`����p�K?���:T�l��2��EF7�lLS��	Q��:MS�ՠ(#Q�K�$���01-A'��,�[3����<**��:�T󾑒�RI�][t����矪� �ǲ��Yẖ�����0"�b�PҘ[B
��p��۩0����`��L�ڜ���a����q�iݧ�8�A8HeB��!�z}u�۶M��Y�'���n�ĊG3X]=�������ͫխV������9??�A��@ɣ�贈a�:��`6F�7�礔�Z-�x�HF��׿2��pH�����ܼy�S��8P|�̉ͯ�ܕ�ٵ�<�����5��2U�XH�8�ÀJ�J���v,�z��(�NZv�T-<�i
Q4"�TVP�{�4lR�湕�|i��B���Klݾ����9�c�峸F��[}l���m�!�2?�Z������>O�V'�$����%G���s�4�sj�H1����{�߻����4j>�c2�P��g��kS��H���TB�|N���1++6+++�޿��8��ѣGsy�;w��.+++�;w�q�
U�6ۖK�L,K2���-s�����t:��y� �s�������n��ƧO]��u�~oĹ��z�a�H��:nN��l[}�˗/�^W�{}nݺ����HŘ�*V��ނ8���k9yZ��:�f�X3��X���F���͛ԫ1/\��n������S~����&�pY\XQ�f���쯔�P���z$���>���5VWW9v�����4}��6�v;�^����
���[ �Y�e�Z�R�Jƣ�h(f���D��&Q����N���S�n�z��F�dIν�]�����v�
A(���x������aܦ��c�����>��D��~�j�Ā�Ԛ��~������f4R�`0ȧ�i#y؀�X��:�Mm�L,JPmԱ��u�$I�����3�>��~�ߔ�����,/]�$/_�,/^�(�(�:��>�}�������[��ߺ,��w�ȗ_{]�˷ORNl�k׾��s��/|��W����߻��z����oO�3=.� �j������<	^{�?j4���������;�v��Y}��B�[�7����"��Z��'������t9�14EG��U�xAzk6ڤ��3��Y�O��6��!�Φ��bW����IF=.tw@�Z��ޫg�O7n�CWpA�0��hFГB���*	�XtΦ�N�1��Cu��8.�`4�L�rt����?K���9-�i�)� ��/Ӈ�\�"?��ʳ��u�u�i��<�@��|�~|Ys�'��5����܇�vv��L�T�6I<y�X�h4Ĕ)�2cF!�����c��2�L�p�ö��5Mϓ<���3�?I7ߓB��گ�$݅O}�i��+iB�WB���F�C����_��ѓF�����ӂ�y�'���:oQ���Mjp��U���d�b��`�w���+���(s=����"s�(vk�y�>.f�`,��F����5-B��M�T4�	C���tiL�=t]G'�tޢ,xރ�f��`�t�g13-�i��Ρξ�Y�z��2PJfY3�����,0����nPj��0m&�noH�H�p�d%�dE	�Wͅ��3m0:��=�A���:�C��&Cj�Z.SV�:�h]�g��vzu�5�_Z�h-��0J���Plڟ��	�qNd�|�2�� ���J�d0��<&��.���3m0Z�R��U=ֈ�z���U�?�ӧOO|�(��̴��n<}E��Sh�kOw ���o��Ǆ�uc�4�03���nY6f��W���M]�Ų,�޽K0����z�k��;-����Lk�l�n���{/��8I��\qt�N�q��Fy߰���}�����!�b�0±l<�x�^�4A0������Z�D��uϗO�.�tv���t���u<K��	S��)e����_�%e�Q�r�3m0�J�P��8U�$�om4zz�$�O��h��`&�z�^�����VY�i���1ד�'M��G�>z��iF��$�j]u]���ݯ�փ\�xTO�i��a��O<7�	A-+�/h�j�}�a�M�,�+�̴�茫�*�C�ȅ�ҒjZ�p1�>���6�l���~��َI�q\�$I҈2*I��*91%O6-��'yB���Q�y�s��he\��|ӆ�7��Tٲ�z���T�CZ,uLf�`tۇ*z�vQ��LL�3�Sa\��|x�DYT�� �i�LGI �j� �0�J/h�E'��q����J~��	�Cв����E�0�8cjҘ��G��?a��>�a����wp���ӥ��Q�!�3}�h����=�Q�$���B�R��Wq]�4��a�ӂ�6-������u�Hk=��6~Mݘ�|�L(�W;�e7�۶��6�b�g�x8���`&�^����j��Xf�,�7��O��&��Sa�(�L[�z�f<s���|tr��I�tY�ƓEc�Ʋ�\��i�B�ϭ�8e��E����3m0��q�����=_d��碈��է���h�vL�x�������L'���T�yQ�l8����H5����N|}���OZ�L��>j��m�Ξ�SD,˿(J�=�a&�ZM���ɢ�#�25t�u�i����I� �^����2�h��8��L�4(t>7�	a8�Uc����� yBM����Q<jd��L��ԽBOÇ�b�_���)NK�&c�78=u{i��#���&���OSY f�`t-GJ���j���H����2	�3m0�b�ia�-֏�c%�����ۍ�m�p��ɈJ�"�4������������Y����+˼x�%���Q�k�A�Z����f���n{�k���s��ܱ�<�k�{��<	f������5N��N�&��8^�z���_=}�4������������f)kmllP��B��/|�Ry̜�H)���R޾}[�axOX&�mq��}�%ʕ���u��666�p��i��o"��:�u�A.�����7���JS�x\�ԕ4�|�0�Vw���2��VJY.BGb[[[�qL��accୌ#3����H����}��$�ˉafN)�Y���E��u����V��S��8{��gΐ�db�]JyU�2Ǖ+W���G���\�t��p���oI)e�2�cY�'~)��R&��������ŋ'�q>5��W�نJ��y    IEND�B`�PK   }Q�TV-&0=  �     jsons/user_defined.json���n�6�_�еH�|�]k��M�(���(*KT�\�߽���wc;��ր/,j�H~C����i퓫d�|�{��P�"I��|ۅ���	�����.�����ǧ�a�}�mV��<k��uS�� ����i�  ���?�wi
s����9#5�k���Bq��B{-4茙��^�����e�;׆u�Mt����E��u}q�P/�I���zxX�n]eO��&�ae�3ٍ�6��Ƃkͷ
ە��� ��bշ�a	��.��^�j�ɬI��f��j��i!�u�U��1`�J6�auz@�cEQ)�s��}�^fU�����jyԀ0 Xk�e��R3NO��?��������R�L�������������/��Q}���5�������ۊ|-��Gm��m^jo,��3��f?�YY7���]L��L�:��9�d(�F �x�$q� ��r���(W�|V+�Xb��*,���-��!�/�ۗ���WfOʿ��W_U�ㄊ�->���jV�^���hL���L΀{��oc�WNS)X��r`�8A��i�DᥧT����� �,��G�'&�Ӂ�p�Q��_RaF4;q?���w��(l4����w���>#�B����b������M=�Y*YQ����@�v�Ȳ� ]:G�ɼ��%�R�|L�D`7g�`� ������j&Si��rq��U���j
��.�Щ��������vv���O�����e�L!�ƚ!åA��<�̗��K������b��R��V�*�h
$���J�Z-�%R�2�c���lJ�30��ET~c�"��2v7w��PK   }Q�TP�d�'  �            ��    cirkitFile.jsonPK   }Q�Ts�7+5J  dK  /           ��(  images/6c71542d-16cb-4630-930f-71c4de5e1144.pngPK   }Q�T��4�� ̻ /           ���r  images/7a4be1c8-201b-41f2-b584-263fc50cb409.pngPK   }Q�T6�0{ { /           ���. images/c51b28eb-c857-4ce7-b81a-d633a3d7e747.pngPK   }Q�T��K� 	� /           ��I� images/cd1eebff-8d4c-4172-8358-6f93b12ef793.pngPK   }Q�T��!�D�  Ԟ  /           ���D images/cf2dd1a8-295d-437f-92b8-7fcc138ae9be.pngPK   }Q�TV-&0=  �             ��r� jsons/user_defined.jsonPK      S  ��   